// Modified by Princeton University on June 9th, 2015
// ========== Copyright Header Begin ==========================================
//
// OpenSPARC T1 Processor File: pc_cmp.v
// Copyright (c) 2006 Sun Microsystems, Inc.  All Rights Reserved.
// DO NOT ALTER OR REMOVE COPYRIGHT NOTICES.
//
// The above named program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public
// License version 2 as published by the Free Software Foundation.
//
// The above named program is distributed in the hope that it will be
// useful, but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
// General Public License for more details.
//
// You should have received a copy of the GNU General Public
// License along with this work; if not, write to the Free Software
// Foundation, Inc., 51 Franklin St, Fifth Floor, Boston, MA 02110-1301, USA.
//
// ========== Copyright Header End ============================================

`include "define.tmp.h"
`include "ifu.tmp.h"

// /home/gl/work/openpiton/piton/verif/env/manycore/devices_ariane.xml
`define GOOD_TRAP_COUNTER 1


 module pc_cmp(/*AUTOARG*/
     // Inputs
     clk,
     rst_l
 );
input clk;
input rst_l;

// trap register

reg [1023:0]   active_thread;
reg [4:0]    thread_status[1023:0];

reg [255:0]   good = '0;
reg [255:0]   done;

reg [31:0]     timeout [1023:0];


reg [63:0]    good_trap[`GOOD_TRAP_COUNTER-1:0];
reg [63:0]    bad_trap [`GOOD_TRAP_COUNTER-1:0];

reg [`GOOD_TRAP_COUNTER-1:0] good_trap_exists;
reg [`GOOD_TRAP_COUNTER-1:0] bad_trap_exists;

reg           dum;
reg           hit_bad = 0;

integer       time_tmp, trap_count;


    reg spc0_inst_done;
    wire [1:0]   spc0_thread_id;
    wire [63:0]      spc0_rtl_pc;
    wire sas_m0;
    reg [63:0] spc0_phy_pc_w;

    

    reg spc1_inst_done;
    wire [1:0]   spc1_thread_id;
    wire [63:0]      spc1_rtl_pc;
    wire sas_m1;
    reg [63:0] spc1_phy_pc_w;

    

    reg spc2_inst_done;
    wire [1:0]   spc2_thread_id;
    wire [63:0]      spc2_rtl_pc;
    wire sas_m2;
    reg [63:0] spc2_phy_pc_w;

    

    reg spc3_inst_done;
    wire [1:0]   spc3_thread_id;
    wire [63:0]      spc3_rtl_pc;
    wire sas_m3;
    reg [63:0] spc3_phy_pc_w;

    

    reg spc4_inst_done;
    wire [1:0]   spc4_thread_id;
    wire [63:0]      spc4_rtl_pc;
    wire sas_m4;
    reg [63:0] spc4_phy_pc_w;

    

    reg spc5_inst_done;
    wire [1:0]   spc5_thread_id;
    wire [63:0]      spc5_rtl_pc;
    wire sas_m5;
    reg [63:0] spc5_phy_pc_w;

    

    reg spc6_inst_done;
    wire [1:0]   spc6_thread_id;
    wire [63:0]      spc6_rtl_pc;
    wire sas_m6;
    reg [63:0] spc6_phy_pc_w;

    

    reg spc7_inst_done;
    wire [1:0]   spc7_thread_id;
    wire [63:0]      spc7_rtl_pc;
    wire sas_m7;
    reg [63:0] spc7_phy_pc_w;

    

    reg spc8_inst_done;
    wire [1:0]   spc8_thread_id;
    wire [63:0]      spc8_rtl_pc;
    wire sas_m8;
    reg [63:0] spc8_phy_pc_w;

    

    reg spc9_inst_done;
    wire [1:0]   spc9_thread_id;
    wire [63:0]      spc9_rtl_pc;
    wire sas_m9;
    reg [63:0] spc9_phy_pc_w;

    

    reg spc10_inst_done;
    wire [1:0]   spc10_thread_id;
    wire [63:0]      spc10_rtl_pc;
    wire sas_m10;
    reg [63:0] spc10_phy_pc_w;

    

    reg spc11_inst_done;
    wire [1:0]   spc11_thread_id;
    wire [63:0]      spc11_rtl_pc;
    wire sas_m11;
    reg [63:0] spc11_phy_pc_w;

    

    reg spc12_inst_done;
    wire [1:0]   spc12_thread_id;
    wire [63:0]      spc12_rtl_pc;
    wire sas_m12;
    reg [63:0] spc12_phy_pc_w;

    

    reg spc13_inst_done;
    wire [1:0]   spc13_thread_id;
    wire [63:0]      spc13_rtl_pc;
    wire sas_m13;
    reg [63:0] spc13_phy_pc_w;

    

    reg spc14_inst_done;
    wire [1:0]   spc14_thread_id;
    wire [63:0]      spc14_rtl_pc;
    wire sas_m14;
    reg [63:0] spc14_phy_pc_w;

    

    reg spc15_inst_done;
    wire [1:0]   spc15_thread_id;
    wire [63:0]      spc15_rtl_pc;
    wire sas_m15;
    reg [63:0] spc15_phy_pc_w;

    

    reg spc16_inst_done;
    wire [1:0]   spc16_thread_id;
    wire [63:0]      spc16_rtl_pc;
    wire sas_m16;
    reg [63:0] spc16_phy_pc_w;

    

    reg spc17_inst_done;
    wire [1:0]   spc17_thread_id;
    wire [63:0]      spc17_rtl_pc;
    wire sas_m17;
    reg [63:0] spc17_phy_pc_w;

    

    reg spc18_inst_done;
    wire [1:0]   spc18_thread_id;
    wire [63:0]      spc18_rtl_pc;
    wire sas_m18;
    reg [63:0] spc18_phy_pc_w;

    

    reg spc19_inst_done;
    wire [1:0]   spc19_thread_id;
    wire [63:0]      spc19_rtl_pc;
    wire sas_m19;
    reg [63:0] spc19_phy_pc_w;

    

    reg spc20_inst_done;
    wire [1:0]   spc20_thread_id;
    wire [63:0]      spc20_rtl_pc;
    wire sas_m20;
    reg [63:0] spc20_phy_pc_w;

    

    reg spc21_inst_done;
    wire [1:0]   spc21_thread_id;
    wire [63:0]      spc21_rtl_pc;
    wire sas_m21;
    reg [63:0] spc21_phy_pc_w;

    

    reg spc22_inst_done;
    wire [1:0]   spc22_thread_id;
    wire [63:0]      spc22_rtl_pc;
    wire sas_m22;
    reg [63:0] spc22_phy_pc_w;

    

    reg spc23_inst_done;
    wire [1:0]   spc23_thread_id;
    wire [63:0]      spc23_rtl_pc;
    wire sas_m23;
    reg [63:0] spc23_phy_pc_w;

    

    reg spc24_inst_done;
    wire [1:0]   spc24_thread_id;
    wire [63:0]      spc24_rtl_pc;
    wire sas_m24;
    reg [63:0] spc24_phy_pc_w;

    

    reg spc25_inst_done;
    wire [1:0]   spc25_thread_id;
    wire [63:0]      spc25_rtl_pc;
    wire sas_m25;
    reg [63:0] spc25_phy_pc_w;

    

    reg spc26_inst_done;
    wire [1:0]   spc26_thread_id;
    wire [63:0]      spc26_rtl_pc;
    wire sas_m26;
    reg [63:0] spc26_phy_pc_w;

    

    reg spc27_inst_done;
    wire [1:0]   spc27_thread_id;
    wire [63:0]      spc27_rtl_pc;
    wire sas_m27;
    reg [63:0] spc27_phy_pc_w;

    

    reg spc28_inst_done;
    wire [1:0]   spc28_thread_id;
    wire [63:0]      spc28_rtl_pc;
    wire sas_m28;
    reg [63:0] spc28_phy_pc_w;

    

    reg spc29_inst_done;
    wire [1:0]   spc29_thread_id;
    wire [63:0]      spc29_rtl_pc;
    wire sas_m29;
    reg [63:0] spc29_phy_pc_w;

    

    reg spc30_inst_done;
    wire [1:0]   spc30_thread_id;
    wire [63:0]      spc30_rtl_pc;
    wire sas_m30;
    reg [63:0] spc30_phy_pc_w;

    

    reg spc31_inst_done;
    wire [1:0]   spc31_thread_id;
    wire [63:0]      spc31_rtl_pc;
    wire sas_m31;
    reg [63:0] spc31_phy_pc_w;

    

    reg spc32_inst_done;
    wire [1:0]   spc32_thread_id;
    wire [63:0]      spc32_rtl_pc;
    wire sas_m32;
    reg [63:0] spc32_phy_pc_w;

    

    reg spc33_inst_done;
    wire [1:0]   spc33_thread_id;
    wire [63:0]      spc33_rtl_pc;
    wire sas_m33;
    reg [63:0] spc33_phy_pc_w;

    

    reg spc34_inst_done;
    wire [1:0]   spc34_thread_id;
    wire [63:0]      spc34_rtl_pc;
    wire sas_m34;
    reg [63:0] spc34_phy_pc_w;

    

    reg spc35_inst_done;
    wire [1:0]   spc35_thread_id;
    wire [63:0]      spc35_rtl_pc;
    wire sas_m35;
    reg [63:0] spc35_phy_pc_w;

    

    reg spc36_inst_done;
    wire [1:0]   spc36_thread_id;
    wire [63:0]      spc36_rtl_pc;
    wire sas_m36;
    reg [63:0] spc36_phy_pc_w;

    

    reg spc37_inst_done;
    wire [1:0]   spc37_thread_id;
    wire [63:0]      spc37_rtl_pc;
    wire sas_m37;
    reg [63:0] spc37_phy_pc_w;

    

    reg spc38_inst_done;
    wire [1:0]   spc38_thread_id;
    wire [63:0]      spc38_rtl_pc;
    wire sas_m38;
    reg [63:0] spc38_phy_pc_w;

    

    reg spc39_inst_done;
    wire [1:0]   spc39_thread_id;
    wire [63:0]      spc39_rtl_pc;
    wire sas_m39;
    reg [63:0] spc39_phy_pc_w;

    

    reg spc40_inst_done;
    wire [1:0]   spc40_thread_id;
    wire [63:0]      spc40_rtl_pc;
    wire sas_m40;
    reg [63:0] spc40_phy_pc_w;

    

    reg spc41_inst_done;
    wire [1:0]   spc41_thread_id;
    wire [63:0]      spc41_rtl_pc;
    wire sas_m41;
    reg [63:0] spc41_phy_pc_w;

    

    reg spc42_inst_done;
    wire [1:0]   spc42_thread_id;
    wire [63:0]      spc42_rtl_pc;
    wire sas_m42;
    reg [63:0] spc42_phy_pc_w;

    

    reg spc43_inst_done;
    wire [1:0]   spc43_thread_id;
    wire [63:0]      spc43_rtl_pc;
    wire sas_m43;
    reg [63:0] spc43_phy_pc_w;

    

    reg spc44_inst_done;
    wire [1:0]   spc44_thread_id;
    wire [63:0]      spc44_rtl_pc;
    wire sas_m44;
    reg [63:0] spc44_phy_pc_w;

    

    reg spc45_inst_done;
    wire [1:0]   spc45_thread_id;
    wire [63:0]      spc45_rtl_pc;
    wire sas_m45;
    reg [63:0] spc45_phy_pc_w;

    

    reg spc46_inst_done;
    wire [1:0]   spc46_thread_id;
    wire [63:0]      spc46_rtl_pc;
    wire sas_m46;
    reg [63:0] spc46_phy_pc_w;

    

    reg spc47_inst_done;
    wire [1:0]   spc47_thread_id;
    wire [63:0]      spc47_rtl_pc;
    wire sas_m47;
    reg [63:0] spc47_phy_pc_w;

    

    reg spc48_inst_done;
    wire [1:0]   spc48_thread_id;
    wire [63:0]      spc48_rtl_pc;
    wire sas_m48;
    reg [63:0] spc48_phy_pc_w;

    

    reg spc49_inst_done;
    wire [1:0]   spc49_thread_id;
    wire [63:0]      spc49_rtl_pc;
    wire sas_m49;
    reg [63:0] spc49_phy_pc_w;

    

    reg spc50_inst_done;
    wire [1:0]   spc50_thread_id;
    wire [63:0]      spc50_rtl_pc;
    wire sas_m50;
    reg [63:0] spc50_phy_pc_w;

    

    reg spc51_inst_done;
    wire [1:0]   spc51_thread_id;
    wire [63:0]      spc51_rtl_pc;
    wire sas_m51;
    reg [63:0] spc51_phy_pc_w;

    

    reg spc52_inst_done;
    wire [1:0]   spc52_thread_id;
    wire [63:0]      spc52_rtl_pc;
    wire sas_m52;
    reg [63:0] spc52_phy_pc_w;

    

    reg spc53_inst_done;
    wire [1:0]   spc53_thread_id;
    wire [63:0]      spc53_rtl_pc;
    wire sas_m53;
    reg [63:0] spc53_phy_pc_w;

    

    reg spc54_inst_done;
    wire [1:0]   spc54_thread_id;
    wire [63:0]      spc54_rtl_pc;
    wire sas_m54;
    reg [63:0] spc54_phy_pc_w;

    

    reg spc55_inst_done;
    wire [1:0]   spc55_thread_id;
    wire [63:0]      spc55_rtl_pc;
    wire sas_m55;
    reg [63:0] spc55_phy_pc_w;

    

    reg spc56_inst_done;
    wire [1:0]   spc56_thread_id;
    wire [63:0]      spc56_rtl_pc;
    wire sas_m56;
    reg [63:0] spc56_phy_pc_w;

    

    reg spc57_inst_done;
    wire [1:0]   spc57_thread_id;
    wire [63:0]      spc57_rtl_pc;
    wire sas_m57;
    reg [63:0] spc57_phy_pc_w;

    

    reg spc58_inst_done;
    wire [1:0]   spc58_thread_id;
    wire [63:0]      spc58_rtl_pc;
    wire sas_m58;
    reg [63:0] spc58_phy_pc_w;

    

    reg spc59_inst_done;
    wire [1:0]   spc59_thread_id;
    wire [63:0]      spc59_rtl_pc;
    wire sas_m59;
    reg [63:0] spc59_phy_pc_w;

    

    reg spc60_inst_done;
    wire [1:0]   spc60_thread_id;
    wire [63:0]      spc60_rtl_pc;
    wire sas_m60;
    reg [63:0] spc60_phy_pc_w;

    

    reg spc61_inst_done;
    wire [1:0]   spc61_thread_id;
    wire [63:0]      spc61_rtl_pc;
    wire sas_m61;
    reg [63:0] spc61_phy_pc_w;

    

    reg spc62_inst_done;
    wire [1:0]   spc62_thread_id;
    wire [63:0]      spc62_rtl_pc;
    wire sas_m62;
    reg [63:0] spc62_phy_pc_w;

    

    reg spc63_inst_done;
    wire [1:0]   spc63_thread_id;
    wire [63:0]      spc63_rtl_pc;
    wire sas_m63;
    reg [63:0] spc63_phy_pc_w;

    

    reg spc64_inst_done;
    wire [1:0]   spc64_thread_id;
    wire [63:0]      spc64_rtl_pc;
    wire sas_m64;
    reg [63:0] spc64_phy_pc_w;

    

    reg spc65_inst_done;
    wire [1:0]   spc65_thread_id;
    wire [63:0]      spc65_rtl_pc;
    wire sas_m65;
    reg [63:0] spc65_phy_pc_w;

    

    reg spc66_inst_done;
    wire [1:0]   spc66_thread_id;
    wire [63:0]      spc66_rtl_pc;
    wire sas_m66;
    reg [63:0] spc66_phy_pc_w;

    

    reg spc67_inst_done;
    wire [1:0]   spc67_thread_id;
    wire [63:0]      spc67_rtl_pc;
    wire sas_m67;
    reg [63:0] spc67_phy_pc_w;

    

    reg spc68_inst_done;
    wire [1:0]   spc68_thread_id;
    wire [63:0]      spc68_rtl_pc;
    wire sas_m68;
    reg [63:0] spc68_phy_pc_w;

    

    reg spc69_inst_done;
    wire [1:0]   spc69_thread_id;
    wire [63:0]      spc69_rtl_pc;
    wire sas_m69;
    reg [63:0] spc69_phy_pc_w;

    

    reg spc70_inst_done;
    wire [1:0]   spc70_thread_id;
    wire [63:0]      spc70_rtl_pc;
    wire sas_m70;
    reg [63:0] spc70_phy_pc_w;

    

    reg spc71_inst_done;
    wire [1:0]   spc71_thread_id;
    wire [63:0]      spc71_rtl_pc;
    wire sas_m71;
    reg [63:0] spc71_phy_pc_w;

    

    reg spc72_inst_done;
    wire [1:0]   spc72_thread_id;
    wire [63:0]      spc72_rtl_pc;
    wire sas_m72;
    reg [63:0] spc72_phy_pc_w;

    

    reg spc73_inst_done;
    wire [1:0]   spc73_thread_id;
    wire [63:0]      spc73_rtl_pc;
    wire sas_m73;
    reg [63:0] spc73_phy_pc_w;

    

    reg spc74_inst_done;
    wire [1:0]   spc74_thread_id;
    wire [63:0]      spc74_rtl_pc;
    wire sas_m74;
    reg [63:0] spc74_phy_pc_w;

    

    reg spc75_inst_done;
    wire [1:0]   spc75_thread_id;
    wire [63:0]      spc75_rtl_pc;
    wire sas_m75;
    reg [63:0] spc75_phy_pc_w;

    

    reg spc76_inst_done;
    wire [1:0]   spc76_thread_id;
    wire [63:0]      spc76_rtl_pc;
    wire sas_m76;
    reg [63:0] spc76_phy_pc_w;

    

    reg spc77_inst_done;
    wire [1:0]   spc77_thread_id;
    wire [63:0]      spc77_rtl_pc;
    wire sas_m77;
    reg [63:0] spc77_phy_pc_w;

    

    reg spc78_inst_done;
    wire [1:0]   spc78_thread_id;
    wire [63:0]      spc78_rtl_pc;
    wire sas_m78;
    reg [63:0] spc78_phy_pc_w;

    

    reg spc79_inst_done;
    wire [1:0]   spc79_thread_id;
    wire [63:0]      spc79_rtl_pc;
    wire sas_m79;
    reg [63:0] spc79_phy_pc_w;

    

    reg spc80_inst_done;
    wire [1:0]   spc80_thread_id;
    wire [63:0]      spc80_rtl_pc;
    wire sas_m80;
    reg [63:0] spc80_phy_pc_w;

    

    reg spc81_inst_done;
    wire [1:0]   spc81_thread_id;
    wire [63:0]      spc81_rtl_pc;
    wire sas_m81;
    reg [63:0] spc81_phy_pc_w;

    

    reg spc82_inst_done;
    wire [1:0]   spc82_thread_id;
    wire [63:0]      spc82_rtl_pc;
    wire sas_m82;
    reg [63:0] spc82_phy_pc_w;

    

    reg spc83_inst_done;
    wire [1:0]   spc83_thread_id;
    wire [63:0]      spc83_rtl_pc;
    wire sas_m83;
    reg [63:0] spc83_phy_pc_w;

    

    reg spc84_inst_done;
    wire [1:0]   spc84_thread_id;
    wire [63:0]      spc84_rtl_pc;
    wire sas_m84;
    reg [63:0] spc84_phy_pc_w;

    

    reg spc85_inst_done;
    wire [1:0]   spc85_thread_id;
    wire [63:0]      spc85_rtl_pc;
    wire sas_m85;
    reg [63:0] spc85_phy_pc_w;

    

    reg spc86_inst_done;
    wire [1:0]   spc86_thread_id;
    wire [63:0]      spc86_rtl_pc;
    wire sas_m86;
    reg [63:0] spc86_phy_pc_w;

    

    reg spc87_inst_done;
    wire [1:0]   spc87_thread_id;
    wire [63:0]      spc87_rtl_pc;
    wire sas_m87;
    reg [63:0] spc87_phy_pc_w;

    

    reg spc88_inst_done;
    wire [1:0]   spc88_thread_id;
    wire [63:0]      spc88_rtl_pc;
    wire sas_m88;
    reg [63:0] spc88_phy_pc_w;

    

    reg spc89_inst_done;
    wire [1:0]   spc89_thread_id;
    wire [63:0]      spc89_rtl_pc;
    wire sas_m89;
    reg [63:0] spc89_phy_pc_w;

    

    reg spc90_inst_done;
    wire [1:0]   spc90_thread_id;
    wire [63:0]      spc90_rtl_pc;
    wire sas_m90;
    reg [63:0] spc90_phy_pc_w;

    

    reg spc91_inst_done;
    wire [1:0]   spc91_thread_id;
    wire [63:0]      spc91_rtl_pc;
    wire sas_m91;
    reg [63:0] spc91_phy_pc_w;

    

    reg spc92_inst_done;
    wire [1:0]   spc92_thread_id;
    wire [63:0]      spc92_rtl_pc;
    wire sas_m92;
    reg [63:0] spc92_phy_pc_w;

    

    reg spc93_inst_done;
    wire [1:0]   spc93_thread_id;
    wire [63:0]      spc93_rtl_pc;
    wire sas_m93;
    reg [63:0] spc93_phy_pc_w;

    

    reg spc94_inst_done;
    wire [1:0]   spc94_thread_id;
    wire [63:0]      spc94_rtl_pc;
    wire sas_m94;
    reg [63:0] spc94_phy_pc_w;

    

    reg spc95_inst_done;
    wire [1:0]   spc95_thread_id;
    wire [63:0]      spc95_rtl_pc;
    wire sas_m95;
    reg [63:0] spc95_phy_pc_w;

    

    reg spc96_inst_done;
    wire [1:0]   spc96_thread_id;
    wire [63:0]      spc96_rtl_pc;
    wire sas_m96;
    reg [63:0] spc96_phy_pc_w;

    

    reg spc97_inst_done;
    wire [1:0]   spc97_thread_id;
    wire [63:0]      spc97_rtl_pc;
    wire sas_m97;
    reg [63:0] spc97_phy_pc_w;

    

    reg spc98_inst_done;
    wire [1:0]   spc98_thread_id;
    wire [63:0]      spc98_rtl_pc;
    wire sas_m98;
    reg [63:0] spc98_phy_pc_w;

    

    reg spc99_inst_done;
    wire [1:0]   spc99_thread_id;
    wire [63:0]      spc99_rtl_pc;
    wire sas_m99;
    reg [63:0] spc99_phy_pc_w;

    

    reg spc100_inst_done;
    wire [1:0]   spc100_thread_id;
    wire [63:0]      spc100_rtl_pc;
    wire sas_m100;
    reg [63:0] spc100_phy_pc_w;

    

    reg spc101_inst_done;
    wire [1:0]   spc101_thread_id;
    wire [63:0]      spc101_rtl_pc;
    wire sas_m101;
    reg [63:0] spc101_phy_pc_w;

    

    reg spc102_inst_done;
    wire [1:0]   spc102_thread_id;
    wire [63:0]      spc102_rtl_pc;
    wire sas_m102;
    reg [63:0] spc102_phy_pc_w;

    

    reg spc103_inst_done;
    wire [1:0]   spc103_thread_id;
    wire [63:0]      spc103_rtl_pc;
    wire sas_m103;
    reg [63:0] spc103_phy_pc_w;

    

    reg spc104_inst_done;
    wire [1:0]   spc104_thread_id;
    wire [63:0]      spc104_rtl_pc;
    wire sas_m104;
    reg [63:0] spc104_phy_pc_w;

    

    reg spc105_inst_done;
    wire [1:0]   spc105_thread_id;
    wire [63:0]      spc105_rtl_pc;
    wire sas_m105;
    reg [63:0] spc105_phy_pc_w;

    

    reg spc106_inst_done;
    wire [1:0]   spc106_thread_id;
    wire [63:0]      spc106_rtl_pc;
    wire sas_m106;
    reg [63:0] spc106_phy_pc_w;

    

    reg spc107_inst_done;
    wire [1:0]   spc107_thread_id;
    wire [63:0]      spc107_rtl_pc;
    wire sas_m107;
    reg [63:0] spc107_phy_pc_w;

    

    reg spc108_inst_done;
    wire [1:0]   spc108_thread_id;
    wire [63:0]      spc108_rtl_pc;
    wire sas_m108;
    reg [63:0] spc108_phy_pc_w;

    

    reg spc109_inst_done;
    wire [1:0]   spc109_thread_id;
    wire [63:0]      spc109_rtl_pc;
    wire sas_m109;
    reg [63:0] spc109_phy_pc_w;

    

    reg spc110_inst_done;
    wire [1:0]   spc110_thread_id;
    wire [63:0]      spc110_rtl_pc;
    wire sas_m110;
    reg [63:0] spc110_phy_pc_w;

    

    reg spc111_inst_done;
    wire [1:0]   spc111_thread_id;
    wire [63:0]      spc111_rtl_pc;
    wire sas_m111;
    reg [63:0] spc111_phy_pc_w;

    

    reg spc112_inst_done;
    wire [1:0]   spc112_thread_id;
    wire [63:0]      spc112_rtl_pc;
    wire sas_m112;
    reg [63:0] spc112_phy_pc_w;

    

    reg spc113_inst_done;
    wire [1:0]   spc113_thread_id;
    wire [63:0]      spc113_rtl_pc;
    wire sas_m113;
    reg [63:0] spc113_phy_pc_w;

    

    reg spc114_inst_done;
    wire [1:0]   spc114_thread_id;
    wire [63:0]      spc114_rtl_pc;
    wire sas_m114;
    reg [63:0] spc114_phy_pc_w;

    

    reg spc115_inst_done;
    wire [1:0]   spc115_thread_id;
    wire [63:0]      spc115_rtl_pc;
    wire sas_m115;
    reg [63:0] spc115_phy_pc_w;

    

    reg spc116_inst_done;
    wire [1:0]   spc116_thread_id;
    wire [63:0]      spc116_rtl_pc;
    wire sas_m116;
    reg [63:0] spc116_phy_pc_w;

    

    reg spc117_inst_done;
    wire [1:0]   spc117_thread_id;
    wire [63:0]      spc117_rtl_pc;
    wire sas_m117;
    reg [63:0] spc117_phy_pc_w;

    

    reg spc118_inst_done;
    wire [1:0]   spc118_thread_id;
    wire [63:0]      spc118_rtl_pc;
    wire sas_m118;
    reg [63:0] spc118_phy_pc_w;

    

    reg spc119_inst_done;
    wire [1:0]   spc119_thread_id;
    wire [63:0]      spc119_rtl_pc;
    wire sas_m119;
    reg [63:0] spc119_phy_pc_w;

    

    reg spc120_inst_done;
    wire [1:0]   spc120_thread_id;
    wire [63:0]      spc120_rtl_pc;
    wire sas_m120;
    reg [63:0] spc120_phy_pc_w;

    

    reg spc121_inst_done;
    wire [1:0]   spc121_thread_id;
    wire [63:0]      spc121_rtl_pc;
    wire sas_m121;
    reg [63:0] spc121_phy_pc_w;

    

    reg spc122_inst_done;
    wire [1:0]   spc122_thread_id;
    wire [63:0]      spc122_rtl_pc;
    wire sas_m122;
    reg [63:0] spc122_phy_pc_w;

    

    reg spc123_inst_done;
    wire [1:0]   spc123_thread_id;
    wire [63:0]      spc123_rtl_pc;
    wire sas_m123;
    reg [63:0] spc123_phy_pc_w;

    

    reg spc124_inst_done;
    wire [1:0]   spc124_thread_id;
    wire [63:0]      spc124_rtl_pc;
    wire sas_m124;
    reg [63:0] spc124_phy_pc_w;

    

    reg spc125_inst_done;
    wire [1:0]   spc125_thread_id;
    wire [63:0]      spc125_rtl_pc;
    wire sas_m125;
    reg [63:0] spc125_phy_pc_w;

    

    reg spc126_inst_done;
    wire [1:0]   spc126_thread_id;
    wire [63:0]      spc126_rtl_pc;
    wire sas_m126;
    reg [63:0] spc126_phy_pc_w;

    

    reg spc127_inst_done;
    wire [1:0]   spc127_thread_id;
    wire [63:0]      spc127_rtl_pc;
    wire sas_m127;
    reg [63:0] spc127_phy_pc_w;

    

    reg spc128_inst_done;
    wire [1:0]   spc128_thread_id;
    wire [63:0]      spc128_rtl_pc;
    wire sas_m128;
    reg [63:0] spc128_phy_pc_w;

    

    reg spc129_inst_done;
    wire [1:0]   spc129_thread_id;
    wire [63:0]      spc129_rtl_pc;
    wire sas_m129;
    reg [63:0] spc129_phy_pc_w;

    

    reg spc130_inst_done;
    wire [1:0]   spc130_thread_id;
    wire [63:0]      spc130_rtl_pc;
    wire sas_m130;
    reg [63:0] spc130_phy_pc_w;

    

    reg spc131_inst_done;
    wire [1:0]   spc131_thread_id;
    wire [63:0]      spc131_rtl_pc;
    wire sas_m131;
    reg [63:0] spc131_phy_pc_w;

    

    reg spc132_inst_done;
    wire [1:0]   spc132_thread_id;
    wire [63:0]      spc132_rtl_pc;
    wire sas_m132;
    reg [63:0] spc132_phy_pc_w;

    

    reg spc133_inst_done;
    wire [1:0]   spc133_thread_id;
    wire [63:0]      spc133_rtl_pc;
    wire sas_m133;
    reg [63:0] spc133_phy_pc_w;

    

    reg spc134_inst_done;
    wire [1:0]   spc134_thread_id;
    wire [63:0]      spc134_rtl_pc;
    wire sas_m134;
    reg [63:0] spc134_phy_pc_w;

    

    reg spc135_inst_done;
    wire [1:0]   spc135_thread_id;
    wire [63:0]      spc135_rtl_pc;
    wire sas_m135;
    reg [63:0] spc135_phy_pc_w;

    

    reg spc136_inst_done;
    wire [1:0]   spc136_thread_id;
    wire [63:0]      spc136_rtl_pc;
    wire sas_m136;
    reg [63:0] spc136_phy_pc_w;

    

    reg spc137_inst_done;
    wire [1:0]   spc137_thread_id;
    wire [63:0]      spc137_rtl_pc;
    wire sas_m137;
    reg [63:0] spc137_phy_pc_w;

    

    reg spc138_inst_done;
    wire [1:0]   spc138_thread_id;
    wire [63:0]      spc138_rtl_pc;
    wire sas_m138;
    reg [63:0] spc138_phy_pc_w;

    

    reg spc139_inst_done;
    wire [1:0]   spc139_thread_id;
    wire [63:0]      spc139_rtl_pc;
    wire sas_m139;
    reg [63:0] spc139_phy_pc_w;

    

    reg spc140_inst_done;
    wire [1:0]   spc140_thread_id;
    wire [63:0]      spc140_rtl_pc;
    wire sas_m140;
    reg [63:0] spc140_phy_pc_w;

    

    reg spc141_inst_done;
    wire [1:0]   spc141_thread_id;
    wire [63:0]      spc141_rtl_pc;
    wire sas_m141;
    reg [63:0] spc141_phy_pc_w;

    

    reg spc142_inst_done;
    wire [1:0]   spc142_thread_id;
    wire [63:0]      spc142_rtl_pc;
    wire sas_m142;
    reg [63:0] spc142_phy_pc_w;

    

    reg spc143_inst_done;
    wire [1:0]   spc143_thread_id;
    wire [63:0]      spc143_rtl_pc;
    wire sas_m143;
    reg [63:0] spc143_phy_pc_w;

    

    reg spc144_inst_done;
    wire [1:0]   spc144_thread_id;
    wire [63:0]      spc144_rtl_pc;
    wire sas_m144;
    reg [63:0] spc144_phy_pc_w;

    

    reg spc145_inst_done;
    wire [1:0]   spc145_thread_id;
    wire [63:0]      spc145_rtl_pc;
    wire sas_m145;
    reg [63:0] spc145_phy_pc_w;

    

    reg spc146_inst_done;
    wire [1:0]   spc146_thread_id;
    wire [63:0]      spc146_rtl_pc;
    wire sas_m146;
    reg [63:0] spc146_phy_pc_w;

    

    reg spc147_inst_done;
    wire [1:0]   spc147_thread_id;
    wire [63:0]      spc147_rtl_pc;
    wire sas_m147;
    reg [63:0] spc147_phy_pc_w;

    

    reg spc148_inst_done;
    wire [1:0]   spc148_thread_id;
    wire [63:0]      spc148_rtl_pc;
    wire sas_m148;
    reg [63:0] spc148_phy_pc_w;

    

    reg spc149_inst_done;
    wire [1:0]   spc149_thread_id;
    wire [63:0]      spc149_rtl_pc;
    wire sas_m149;
    reg [63:0] spc149_phy_pc_w;

    

    reg spc150_inst_done;
    wire [1:0]   spc150_thread_id;
    wire [63:0]      spc150_rtl_pc;
    wire sas_m150;
    reg [63:0] spc150_phy_pc_w;

    

    reg spc151_inst_done;
    wire [1:0]   spc151_thread_id;
    wire [63:0]      spc151_rtl_pc;
    wire sas_m151;
    reg [63:0] spc151_phy_pc_w;

    

    reg spc152_inst_done;
    wire [1:0]   spc152_thread_id;
    wire [63:0]      spc152_rtl_pc;
    wire sas_m152;
    reg [63:0] spc152_phy_pc_w;

    

    reg spc153_inst_done;
    wire [1:0]   spc153_thread_id;
    wire [63:0]      spc153_rtl_pc;
    wire sas_m153;
    reg [63:0] spc153_phy_pc_w;

    

    reg spc154_inst_done;
    wire [1:0]   spc154_thread_id;
    wire [63:0]      spc154_rtl_pc;
    wire sas_m154;
    reg [63:0] spc154_phy_pc_w;

    

    reg spc155_inst_done;
    wire [1:0]   spc155_thread_id;
    wire [63:0]      spc155_rtl_pc;
    wire sas_m155;
    reg [63:0] spc155_phy_pc_w;

    

    reg spc156_inst_done;
    wire [1:0]   spc156_thread_id;
    wire [63:0]      spc156_rtl_pc;
    wire sas_m156;
    reg [63:0] spc156_phy_pc_w;

    

    reg spc157_inst_done;
    wire [1:0]   spc157_thread_id;
    wire [63:0]      spc157_rtl_pc;
    wire sas_m157;
    reg [63:0] spc157_phy_pc_w;

    

    reg spc158_inst_done;
    wire [1:0]   spc158_thread_id;
    wire [63:0]      spc158_rtl_pc;
    wire sas_m158;
    reg [63:0] spc158_phy_pc_w;

    

    reg spc159_inst_done;
    wire [1:0]   spc159_thread_id;
    wire [63:0]      spc159_rtl_pc;
    wire sas_m159;
    reg [63:0] spc159_phy_pc_w;

    

    reg spc160_inst_done;
    wire [1:0]   spc160_thread_id;
    wire [63:0]      spc160_rtl_pc;
    wire sas_m160;
    reg [63:0] spc160_phy_pc_w;

    

    reg spc161_inst_done;
    wire [1:0]   spc161_thread_id;
    wire [63:0]      spc161_rtl_pc;
    wire sas_m161;
    reg [63:0] spc161_phy_pc_w;

    

    reg spc162_inst_done;
    wire [1:0]   spc162_thread_id;
    wire [63:0]      spc162_rtl_pc;
    wire sas_m162;
    reg [63:0] spc162_phy_pc_w;

    

    reg spc163_inst_done;
    wire [1:0]   spc163_thread_id;
    wire [63:0]      spc163_rtl_pc;
    wire sas_m163;
    reg [63:0] spc163_phy_pc_w;

    

    reg spc164_inst_done;
    wire [1:0]   spc164_thread_id;
    wire [63:0]      spc164_rtl_pc;
    wire sas_m164;
    reg [63:0] spc164_phy_pc_w;

    

    reg spc165_inst_done;
    wire [1:0]   spc165_thread_id;
    wire [63:0]      spc165_rtl_pc;
    wire sas_m165;
    reg [63:0] spc165_phy_pc_w;

    

    reg spc166_inst_done;
    wire [1:0]   spc166_thread_id;
    wire [63:0]      spc166_rtl_pc;
    wire sas_m166;
    reg [63:0] spc166_phy_pc_w;

    

    reg spc167_inst_done;
    wire [1:0]   spc167_thread_id;
    wire [63:0]      spc167_rtl_pc;
    wire sas_m167;
    reg [63:0] spc167_phy_pc_w;

    

    reg spc168_inst_done;
    wire [1:0]   spc168_thread_id;
    wire [63:0]      spc168_rtl_pc;
    wire sas_m168;
    reg [63:0] spc168_phy_pc_w;

    

    reg spc169_inst_done;
    wire [1:0]   spc169_thread_id;
    wire [63:0]      spc169_rtl_pc;
    wire sas_m169;
    reg [63:0] spc169_phy_pc_w;

    

    reg spc170_inst_done;
    wire [1:0]   spc170_thread_id;
    wire [63:0]      spc170_rtl_pc;
    wire sas_m170;
    reg [63:0] spc170_phy_pc_w;

    

    reg spc171_inst_done;
    wire [1:0]   spc171_thread_id;
    wire [63:0]      spc171_rtl_pc;
    wire sas_m171;
    reg [63:0] spc171_phy_pc_w;

    

    reg spc172_inst_done;
    wire [1:0]   spc172_thread_id;
    wire [63:0]      spc172_rtl_pc;
    wire sas_m172;
    reg [63:0] spc172_phy_pc_w;

    

    reg spc173_inst_done;
    wire [1:0]   spc173_thread_id;
    wire [63:0]      spc173_rtl_pc;
    wire sas_m173;
    reg [63:0] spc173_phy_pc_w;

    

    reg spc174_inst_done;
    wire [1:0]   spc174_thread_id;
    wire [63:0]      spc174_rtl_pc;
    wire sas_m174;
    reg [63:0] spc174_phy_pc_w;

    

    reg spc175_inst_done;
    wire [1:0]   spc175_thread_id;
    wire [63:0]      spc175_rtl_pc;
    wire sas_m175;
    reg [63:0] spc175_phy_pc_w;

    

    reg spc176_inst_done;
    wire [1:0]   spc176_thread_id;
    wire [63:0]      spc176_rtl_pc;
    wire sas_m176;
    reg [63:0] spc176_phy_pc_w;

    

    reg spc177_inst_done;
    wire [1:0]   spc177_thread_id;
    wire [63:0]      spc177_rtl_pc;
    wire sas_m177;
    reg [63:0] spc177_phy_pc_w;

    

    reg spc178_inst_done;
    wire [1:0]   spc178_thread_id;
    wire [63:0]      spc178_rtl_pc;
    wire sas_m178;
    reg [63:0] spc178_phy_pc_w;

    

    reg spc179_inst_done;
    wire [1:0]   spc179_thread_id;
    wire [63:0]      spc179_rtl_pc;
    wire sas_m179;
    reg [63:0] spc179_phy_pc_w;

    

    reg spc180_inst_done;
    wire [1:0]   spc180_thread_id;
    wire [63:0]      spc180_rtl_pc;
    wire sas_m180;
    reg [63:0] spc180_phy_pc_w;

    

    reg spc181_inst_done;
    wire [1:0]   spc181_thread_id;
    wire [63:0]      spc181_rtl_pc;
    wire sas_m181;
    reg [63:0] spc181_phy_pc_w;

    

    reg spc182_inst_done;
    wire [1:0]   spc182_thread_id;
    wire [63:0]      spc182_rtl_pc;
    wire sas_m182;
    reg [63:0] spc182_phy_pc_w;

    

    reg spc183_inst_done;
    wire [1:0]   spc183_thread_id;
    wire [63:0]      spc183_rtl_pc;
    wire sas_m183;
    reg [63:0] spc183_phy_pc_w;

    

    reg spc184_inst_done;
    wire [1:0]   spc184_thread_id;
    wire [63:0]      spc184_rtl_pc;
    wire sas_m184;
    reg [63:0] spc184_phy_pc_w;

    

    reg spc185_inst_done;
    wire [1:0]   spc185_thread_id;
    wire [63:0]      spc185_rtl_pc;
    wire sas_m185;
    reg [63:0] spc185_phy_pc_w;

    

    reg spc186_inst_done;
    wire [1:0]   spc186_thread_id;
    wire [63:0]      spc186_rtl_pc;
    wire sas_m186;
    reg [63:0] spc186_phy_pc_w;

    

    reg spc187_inst_done;
    wire [1:0]   spc187_thread_id;
    wire [63:0]      spc187_rtl_pc;
    wire sas_m187;
    reg [63:0] spc187_phy_pc_w;

    

    reg spc188_inst_done;
    wire [1:0]   spc188_thread_id;
    wire [63:0]      spc188_rtl_pc;
    wire sas_m188;
    reg [63:0] spc188_phy_pc_w;

    

    reg spc189_inst_done;
    wire [1:0]   spc189_thread_id;
    wire [63:0]      spc189_rtl_pc;
    wire sas_m189;
    reg [63:0] spc189_phy_pc_w;

    

    reg spc190_inst_done;
    wire [1:0]   spc190_thread_id;
    wire [63:0]      spc190_rtl_pc;
    wire sas_m190;
    reg [63:0] spc190_phy_pc_w;

    

    reg spc191_inst_done;
    wire [1:0]   spc191_thread_id;
    wire [63:0]      spc191_rtl_pc;
    wire sas_m191;
    reg [63:0] spc191_phy_pc_w;

    

    reg spc192_inst_done;
    wire [1:0]   spc192_thread_id;
    wire [63:0]      spc192_rtl_pc;
    wire sas_m192;
    reg [63:0] spc192_phy_pc_w;

    

    reg spc193_inst_done;
    wire [1:0]   spc193_thread_id;
    wire [63:0]      spc193_rtl_pc;
    wire sas_m193;
    reg [63:0] spc193_phy_pc_w;

    

    reg spc194_inst_done;
    wire [1:0]   spc194_thread_id;
    wire [63:0]      spc194_rtl_pc;
    wire sas_m194;
    reg [63:0] spc194_phy_pc_w;

    

    reg spc195_inst_done;
    wire [1:0]   spc195_thread_id;
    wire [63:0]      spc195_rtl_pc;
    wire sas_m195;
    reg [63:0] spc195_phy_pc_w;

    

    reg spc196_inst_done;
    wire [1:0]   spc196_thread_id;
    wire [63:0]      spc196_rtl_pc;
    wire sas_m196;
    reg [63:0] spc196_phy_pc_w;

    

    reg spc197_inst_done;
    wire [1:0]   spc197_thread_id;
    wire [63:0]      spc197_rtl_pc;
    wire sas_m197;
    reg [63:0] spc197_phy_pc_w;

    

    reg spc198_inst_done;
    wire [1:0]   spc198_thread_id;
    wire [63:0]      spc198_rtl_pc;
    wire sas_m198;
    reg [63:0] spc198_phy_pc_w;

    

    reg spc199_inst_done;
    wire [1:0]   spc199_thread_id;
    wire [63:0]      spc199_rtl_pc;
    wire sas_m199;
    reg [63:0] spc199_phy_pc_w;

    

    reg spc200_inst_done;
    wire [1:0]   spc200_thread_id;
    wire [63:0]      spc200_rtl_pc;
    wire sas_m200;
    reg [63:0] spc200_phy_pc_w;

    

    reg spc201_inst_done;
    wire [1:0]   spc201_thread_id;
    wire [63:0]      spc201_rtl_pc;
    wire sas_m201;
    reg [63:0] spc201_phy_pc_w;

    

    reg spc202_inst_done;
    wire [1:0]   spc202_thread_id;
    wire [63:0]      spc202_rtl_pc;
    wire sas_m202;
    reg [63:0] spc202_phy_pc_w;

    

    reg spc203_inst_done;
    wire [1:0]   spc203_thread_id;
    wire [63:0]      spc203_rtl_pc;
    wire sas_m203;
    reg [63:0] spc203_phy_pc_w;

    

    reg spc204_inst_done;
    wire [1:0]   spc204_thread_id;
    wire [63:0]      spc204_rtl_pc;
    wire sas_m204;
    reg [63:0] spc204_phy_pc_w;

    

    reg spc205_inst_done;
    wire [1:0]   spc205_thread_id;
    wire [63:0]      spc205_rtl_pc;
    wire sas_m205;
    reg [63:0] spc205_phy_pc_w;

    

    reg spc206_inst_done;
    wire [1:0]   spc206_thread_id;
    wire [63:0]      spc206_rtl_pc;
    wire sas_m206;
    reg [63:0] spc206_phy_pc_w;

    

    reg spc207_inst_done;
    wire [1:0]   spc207_thread_id;
    wire [63:0]      spc207_rtl_pc;
    wire sas_m207;
    reg [63:0] spc207_phy_pc_w;

    

    reg spc208_inst_done;
    wire [1:0]   spc208_thread_id;
    wire [63:0]      spc208_rtl_pc;
    wire sas_m208;
    reg [63:0] spc208_phy_pc_w;

    

    reg spc209_inst_done;
    wire [1:0]   spc209_thread_id;
    wire [63:0]      spc209_rtl_pc;
    wire sas_m209;
    reg [63:0] spc209_phy_pc_w;

    

    reg spc210_inst_done;
    wire [1:0]   spc210_thread_id;
    wire [63:0]      spc210_rtl_pc;
    wire sas_m210;
    reg [63:0] spc210_phy_pc_w;

    

    reg spc211_inst_done;
    wire [1:0]   spc211_thread_id;
    wire [63:0]      spc211_rtl_pc;
    wire sas_m211;
    reg [63:0] spc211_phy_pc_w;

    

    reg spc212_inst_done;
    wire [1:0]   spc212_thread_id;
    wire [63:0]      spc212_rtl_pc;
    wire sas_m212;
    reg [63:0] spc212_phy_pc_w;

    

    reg spc213_inst_done;
    wire [1:0]   spc213_thread_id;
    wire [63:0]      spc213_rtl_pc;
    wire sas_m213;
    reg [63:0] spc213_phy_pc_w;

    

    reg spc214_inst_done;
    wire [1:0]   spc214_thread_id;
    wire [63:0]      spc214_rtl_pc;
    wire sas_m214;
    reg [63:0] spc214_phy_pc_w;

    

    reg spc215_inst_done;
    wire [1:0]   spc215_thread_id;
    wire [63:0]      spc215_rtl_pc;
    wire sas_m215;
    reg [63:0] spc215_phy_pc_w;

    

    reg spc216_inst_done;
    wire [1:0]   spc216_thread_id;
    wire [63:0]      spc216_rtl_pc;
    wire sas_m216;
    reg [63:0] spc216_phy_pc_w;

    

    reg spc217_inst_done;
    wire [1:0]   spc217_thread_id;
    wire [63:0]      spc217_rtl_pc;
    wire sas_m217;
    reg [63:0] spc217_phy_pc_w;

    

    reg spc218_inst_done;
    wire [1:0]   spc218_thread_id;
    wire [63:0]      spc218_rtl_pc;
    wire sas_m218;
    reg [63:0] spc218_phy_pc_w;

    

    reg spc219_inst_done;
    wire [1:0]   spc219_thread_id;
    wire [63:0]      spc219_rtl_pc;
    wire sas_m219;
    reg [63:0] spc219_phy_pc_w;

    

    reg spc220_inst_done;
    wire [1:0]   spc220_thread_id;
    wire [63:0]      spc220_rtl_pc;
    wire sas_m220;
    reg [63:0] spc220_phy_pc_w;

    

    reg spc221_inst_done;
    wire [1:0]   spc221_thread_id;
    wire [63:0]      spc221_rtl_pc;
    wire sas_m221;
    reg [63:0] spc221_phy_pc_w;

    

    reg spc222_inst_done;
    wire [1:0]   spc222_thread_id;
    wire [63:0]      spc222_rtl_pc;
    wire sas_m222;
    reg [63:0] spc222_phy_pc_w;

    

    reg spc223_inst_done;
    wire [1:0]   spc223_thread_id;
    wire [63:0]      spc223_rtl_pc;
    wire sas_m223;
    reg [63:0] spc223_phy_pc_w;

    

    reg spc224_inst_done;
    wire [1:0]   spc224_thread_id;
    wire [63:0]      spc224_rtl_pc;
    wire sas_m224;
    reg [63:0] spc224_phy_pc_w;

    

    reg spc225_inst_done;
    wire [1:0]   spc225_thread_id;
    wire [63:0]      spc225_rtl_pc;
    wire sas_m225;
    reg [63:0] spc225_phy_pc_w;

    

    reg spc226_inst_done;
    wire [1:0]   spc226_thread_id;
    wire [63:0]      spc226_rtl_pc;
    wire sas_m226;
    reg [63:0] spc226_phy_pc_w;

    

    reg spc227_inst_done;
    wire [1:0]   spc227_thread_id;
    wire [63:0]      spc227_rtl_pc;
    wire sas_m227;
    reg [63:0] spc227_phy_pc_w;

    

    reg spc228_inst_done;
    wire [1:0]   spc228_thread_id;
    wire [63:0]      spc228_rtl_pc;
    wire sas_m228;
    reg [63:0] spc228_phy_pc_w;

    

    reg spc229_inst_done;
    wire [1:0]   spc229_thread_id;
    wire [63:0]      spc229_rtl_pc;
    wire sas_m229;
    reg [63:0] spc229_phy_pc_w;

    

    reg spc230_inst_done;
    wire [1:0]   spc230_thread_id;
    wire [63:0]      spc230_rtl_pc;
    wire sas_m230;
    reg [63:0] spc230_phy_pc_w;

    

    reg spc231_inst_done;
    wire [1:0]   spc231_thread_id;
    wire [63:0]      spc231_rtl_pc;
    wire sas_m231;
    reg [63:0] spc231_phy_pc_w;

    

    reg spc232_inst_done;
    wire [1:0]   spc232_thread_id;
    wire [63:0]      spc232_rtl_pc;
    wire sas_m232;
    reg [63:0] spc232_phy_pc_w;

    

    reg spc233_inst_done;
    wire [1:0]   spc233_thread_id;
    wire [63:0]      spc233_rtl_pc;
    wire sas_m233;
    reg [63:0] spc233_phy_pc_w;

    

    reg spc234_inst_done;
    wire [1:0]   spc234_thread_id;
    wire [63:0]      spc234_rtl_pc;
    wire sas_m234;
    reg [63:0] spc234_phy_pc_w;

    

    reg spc235_inst_done;
    wire [1:0]   spc235_thread_id;
    wire [63:0]      spc235_rtl_pc;
    wire sas_m235;
    reg [63:0] spc235_phy_pc_w;

    

    reg spc236_inst_done;
    wire [1:0]   spc236_thread_id;
    wire [63:0]      spc236_rtl_pc;
    wire sas_m236;
    reg [63:0] spc236_phy_pc_w;

    

    reg spc237_inst_done;
    wire [1:0]   spc237_thread_id;
    wire [63:0]      spc237_rtl_pc;
    wire sas_m237;
    reg [63:0] spc237_phy_pc_w;

    

    reg spc238_inst_done;
    wire [1:0]   spc238_thread_id;
    wire [63:0]      spc238_rtl_pc;
    wire sas_m238;
    reg [63:0] spc238_phy_pc_w;

    

    reg spc239_inst_done;
    wire [1:0]   spc239_thread_id;
    wire [63:0]      spc239_rtl_pc;
    wire sas_m239;
    reg [63:0] spc239_phy_pc_w;

    

    reg spc240_inst_done;
    wire [1:0]   spc240_thread_id;
    wire [63:0]      spc240_rtl_pc;
    wire sas_m240;
    reg [63:0] spc240_phy_pc_w;

    

    reg spc241_inst_done;
    wire [1:0]   spc241_thread_id;
    wire [63:0]      spc241_rtl_pc;
    wire sas_m241;
    reg [63:0] spc241_phy_pc_w;

    

    reg spc242_inst_done;
    wire [1:0]   spc242_thread_id;
    wire [63:0]      spc242_rtl_pc;
    wire sas_m242;
    reg [63:0] spc242_phy_pc_w;

    

    reg spc243_inst_done;
    wire [1:0]   spc243_thread_id;
    wire [63:0]      spc243_rtl_pc;
    wire sas_m243;
    reg [63:0] spc243_phy_pc_w;

    

    reg spc244_inst_done;
    wire [1:0]   spc244_thread_id;
    wire [63:0]      spc244_rtl_pc;
    wire sas_m244;
    reg [63:0] spc244_phy_pc_w;

    

    reg spc245_inst_done;
    wire [1:0]   spc245_thread_id;
    wire [63:0]      spc245_rtl_pc;
    wire sas_m245;
    reg [63:0] spc245_phy_pc_w;

    

    reg spc246_inst_done;
    wire [1:0]   spc246_thread_id;
    wire [63:0]      spc246_rtl_pc;
    wire sas_m246;
    reg [63:0] spc246_phy_pc_w;

    

    reg spc247_inst_done;
    wire [1:0]   spc247_thread_id;
    wire [63:0]      spc247_rtl_pc;
    wire sas_m247;
    reg [63:0] spc247_phy_pc_w;

    

    reg spc248_inst_done;
    wire [1:0]   spc248_thread_id;
    wire [63:0]      spc248_rtl_pc;
    wire sas_m248;
    reg [63:0] spc248_phy_pc_w;

    

    reg spc249_inst_done;
    wire [1:0]   spc249_thread_id;
    wire [63:0]      spc249_rtl_pc;
    wire sas_m249;
    reg [63:0] spc249_phy_pc_w;

    

    reg spc250_inst_done;
    wire [1:0]   spc250_thread_id;
    wire [63:0]      spc250_rtl_pc;
    wire sas_m250;
    reg [63:0] spc250_phy_pc_w;

    

    reg spc251_inst_done;
    wire [1:0]   spc251_thread_id;
    wire [63:0]      spc251_rtl_pc;
    wire sas_m251;
    reg [63:0] spc251_phy_pc_w;

    

    reg spc252_inst_done;
    wire [1:0]   spc252_thread_id;
    wire [63:0]      spc252_rtl_pc;
    wire sas_m252;
    reg [63:0] spc252_phy_pc_w;

    

    reg spc253_inst_done;
    wire [1:0]   spc253_thread_id;
    wire [63:0]      spc253_rtl_pc;
    wire sas_m253;
    reg [63:0] spc253_phy_pc_w;

    

    reg spc254_inst_done;
    wire [1:0]   spc254_thread_id;
    wire [63:0]      spc254_rtl_pc;
    wire sas_m254;
    reg [63:0] spc254_phy_pc_w;

    

    reg spc255_inst_done;
    wire [1:0]   spc255_thread_id;
    wire [63:0]      spc255_rtl_pc;
    wire sas_m255;
    reg [63:0] spc255_phy_pc_w;

    


integer      good_trap_count;
integer      bad_trap_count;
reg         local_diag_done;

//use this for the second reset.
initial begin
    local_diag_done = 0;

    good_trap_exists = {`GOOD_TRAP_COUNTER{1'b0}};
    bad_trap_exists = {`GOOD_TRAP_COUNTER{1'b0}};
end
//-----------------------------------------------------------

`ifdef INCLUDE_SAS_TASKS
task get_thread_status;
    begin
    thread_status[0] = `IFUPATH0.swl.thr0_state;
thread_status[1] = `IFUPATH0.swl.thr1_state;
thread_status[2] = `IFUPATH0.swl.thr2_state;
thread_status[3] = `IFUPATH0.swl.thr3_state;
thread_status[4] = `IFUPATH1.swl.thr0_state;
thread_status[5] = `IFUPATH1.swl.thr1_state;
thread_status[6] = `IFUPATH1.swl.thr2_state;
thread_status[7] = `IFUPATH1.swl.thr3_state;
thread_status[8] = `IFUPATH2.swl.thr0_state;
thread_status[9] = `IFUPATH2.swl.thr1_state;
thread_status[10] = `IFUPATH2.swl.thr2_state;
thread_status[11] = `IFUPATH2.swl.thr3_state;
thread_status[12] = `IFUPATH3.swl.thr0_state;
thread_status[13] = `IFUPATH3.swl.thr1_state;
thread_status[14] = `IFUPATH3.swl.thr2_state;
thread_status[15] = `IFUPATH3.swl.thr3_state;
thread_status[16] = `IFUPATH4.swl.thr0_state;
thread_status[17] = `IFUPATH4.swl.thr1_state;
thread_status[18] = `IFUPATH4.swl.thr2_state;
thread_status[19] = `IFUPATH4.swl.thr3_state;
thread_status[20] = `IFUPATH5.swl.thr0_state;
thread_status[21] = `IFUPATH5.swl.thr1_state;
thread_status[22] = `IFUPATH5.swl.thr2_state;
thread_status[23] = `IFUPATH5.swl.thr3_state;
thread_status[24] = `IFUPATH6.swl.thr0_state;
thread_status[25] = `IFUPATH6.swl.thr1_state;
thread_status[26] = `IFUPATH6.swl.thr2_state;
thread_status[27] = `IFUPATH6.swl.thr3_state;
thread_status[28] = `IFUPATH7.swl.thr0_state;
thread_status[29] = `IFUPATH7.swl.thr1_state;
thread_status[30] = `IFUPATH7.swl.thr2_state;
thread_status[31] = `IFUPATH7.swl.thr3_state;
thread_status[32] = `IFUPATH8.swl.thr0_state;
thread_status[33] = `IFUPATH8.swl.thr1_state;
thread_status[34] = `IFUPATH8.swl.thr2_state;
thread_status[35] = `IFUPATH8.swl.thr3_state;
thread_status[36] = `IFUPATH9.swl.thr0_state;
thread_status[37] = `IFUPATH9.swl.thr1_state;
thread_status[38] = `IFUPATH9.swl.thr2_state;
thread_status[39] = `IFUPATH9.swl.thr3_state;
thread_status[40] = `IFUPATH10.swl.thr0_state;
thread_status[41] = `IFUPATH10.swl.thr1_state;
thread_status[42] = `IFUPATH10.swl.thr2_state;
thread_status[43] = `IFUPATH10.swl.thr3_state;
thread_status[44] = `IFUPATH11.swl.thr0_state;
thread_status[45] = `IFUPATH11.swl.thr1_state;
thread_status[46] = `IFUPATH11.swl.thr2_state;
thread_status[47] = `IFUPATH11.swl.thr3_state;
thread_status[48] = `IFUPATH12.swl.thr0_state;
thread_status[49] = `IFUPATH12.swl.thr1_state;
thread_status[50] = `IFUPATH12.swl.thr2_state;
thread_status[51] = `IFUPATH12.swl.thr3_state;
thread_status[52] = `IFUPATH13.swl.thr0_state;
thread_status[53] = `IFUPATH13.swl.thr1_state;
thread_status[54] = `IFUPATH13.swl.thr2_state;
thread_status[55] = `IFUPATH13.swl.thr3_state;
thread_status[56] = `IFUPATH14.swl.thr0_state;
thread_status[57] = `IFUPATH14.swl.thr1_state;
thread_status[58] = `IFUPATH14.swl.thr2_state;
thread_status[59] = `IFUPATH14.swl.thr3_state;
thread_status[60] = `IFUPATH15.swl.thr0_state;
thread_status[61] = `IFUPATH15.swl.thr1_state;
thread_status[62] = `IFUPATH15.swl.thr2_state;
thread_status[63] = `IFUPATH15.swl.thr3_state;
thread_status[64] = `IFUPATH16.swl.thr0_state;
thread_status[65] = `IFUPATH16.swl.thr1_state;
thread_status[66] = `IFUPATH16.swl.thr2_state;
thread_status[67] = `IFUPATH16.swl.thr3_state;
thread_status[68] = `IFUPATH17.swl.thr0_state;
thread_status[69] = `IFUPATH17.swl.thr1_state;
thread_status[70] = `IFUPATH17.swl.thr2_state;
thread_status[71] = `IFUPATH17.swl.thr3_state;
thread_status[72] = `IFUPATH18.swl.thr0_state;
thread_status[73] = `IFUPATH18.swl.thr1_state;
thread_status[74] = `IFUPATH18.swl.thr2_state;
thread_status[75] = `IFUPATH18.swl.thr3_state;
thread_status[76] = `IFUPATH19.swl.thr0_state;
thread_status[77] = `IFUPATH19.swl.thr1_state;
thread_status[78] = `IFUPATH19.swl.thr2_state;
thread_status[79] = `IFUPATH19.swl.thr3_state;
thread_status[80] = `IFUPATH20.swl.thr0_state;
thread_status[81] = `IFUPATH20.swl.thr1_state;
thread_status[82] = `IFUPATH20.swl.thr2_state;
thread_status[83] = `IFUPATH20.swl.thr3_state;
thread_status[84] = `IFUPATH21.swl.thr0_state;
thread_status[85] = `IFUPATH21.swl.thr1_state;
thread_status[86] = `IFUPATH21.swl.thr2_state;
thread_status[87] = `IFUPATH21.swl.thr3_state;
thread_status[88] = `IFUPATH22.swl.thr0_state;
thread_status[89] = `IFUPATH22.swl.thr1_state;
thread_status[90] = `IFUPATH22.swl.thr2_state;
thread_status[91] = `IFUPATH22.swl.thr3_state;
thread_status[92] = `IFUPATH23.swl.thr0_state;
thread_status[93] = `IFUPATH23.swl.thr1_state;
thread_status[94] = `IFUPATH23.swl.thr2_state;
thread_status[95] = `IFUPATH23.swl.thr3_state;
thread_status[96] = `IFUPATH24.swl.thr0_state;
thread_status[97] = `IFUPATH24.swl.thr1_state;
thread_status[98] = `IFUPATH24.swl.thr2_state;
thread_status[99] = `IFUPATH24.swl.thr3_state;
thread_status[100] = `IFUPATH25.swl.thr0_state;
thread_status[101] = `IFUPATH25.swl.thr1_state;
thread_status[102] = `IFUPATH25.swl.thr2_state;
thread_status[103] = `IFUPATH25.swl.thr3_state;
thread_status[104] = `IFUPATH26.swl.thr0_state;
thread_status[105] = `IFUPATH26.swl.thr1_state;
thread_status[106] = `IFUPATH26.swl.thr2_state;
thread_status[107] = `IFUPATH26.swl.thr3_state;
thread_status[108] = `IFUPATH27.swl.thr0_state;
thread_status[109] = `IFUPATH27.swl.thr1_state;
thread_status[110] = `IFUPATH27.swl.thr2_state;
thread_status[111] = `IFUPATH27.swl.thr3_state;
thread_status[112] = `IFUPATH28.swl.thr0_state;
thread_status[113] = `IFUPATH28.swl.thr1_state;
thread_status[114] = `IFUPATH28.swl.thr2_state;
thread_status[115] = `IFUPATH28.swl.thr3_state;
thread_status[116] = `IFUPATH29.swl.thr0_state;
thread_status[117] = `IFUPATH29.swl.thr1_state;
thread_status[118] = `IFUPATH29.swl.thr2_state;
thread_status[119] = `IFUPATH29.swl.thr3_state;
thread_status[120] = `IFUPATH30.swl.thr0_state;
thread_status[121] = `IFUPATH30.swl.thr1_state;
thread_status[122] = `IFUPATH30.swl.thr2_state;
thread_status[123] = `IFUPATH30.swl.thr3_state;
thread_status[124] = `IFUPATH31.swl.thr0_state;
thread_status[125] = `IFUPATH31.swl.thr1_state;
thread_status[126] = `IFUPATH31.swl.thr2_state;
thread_status[127] = `IFUPATH31.swl.thr3_state;
thread_status[128] = `IFUPATH32.swl.thr0_state;
thread_status[129] = `IFUPATH32.swl.thr1_state;
thread_status[130] = `IFUPATH32.swl.thr2_state;
thread_status[131] = `IFUPATH32.swl.thr3_state;
thread_status[132] = `IFUPATH33.swl.thr0_state;
thread_status[133] = `IFUPATH33.swl.thr1_state;
thread_status[134] = `IFUPATH33.swl.thr2_state;
thread_status[135] = `IFUPATH33.swl.thr3_state;
thread_status[136] = `IFUPATH34.swl.thr0_state;
thread_status[137] = `IFUPATH34.swl.thr1_state;
thread_status[138] = `IFUPATH34.swl.thr2_state;
thread_status[139] = `IFUPATH34.swl.thr3_state;
thread_status[140] = `IFUPATH35.swl.thr0_state;
thread_status[141] = `IFUPATH35.swl.thr1_state;
thread_status[142] = `IFUPATH35.swl.thr2_state;
thread_status[143] = `IFUPATH35.swl.thr3_state;
thread_status[144] = `IFUPATH36.swl.thr0_state;
thread_status[145] = `IFUPATH36.swl.thr1_state;
thread_status[146] = `IFUPATH36.swl.thr2_state;
thread_status[147] = `IFUPATH36.swl.thr3_state;
thread_status[148] = `IFUPATH37.swl.thr0_state;
thread_status[149] = `IFUPATH37.swl.thr1_state;
thread_status[150] = `IFUPATH37.swl.thr2_state;
thread_status[151] = `IFUPATH37.swl.thr3_state;
thread_status[152] = `IFUPATH38.swl.thr0_state;
thread_status[153] = `IFUPATH38.swl.thr1_state;
thread_status[154] = `IFUPATH38.swl.thr2_state;
thread_status[155] = `IFUPATH38.swl.thr3_state;
thread_status[156] = `IFUPATH39.swl.thr0_state;
thread_status[157] = `IFUPATH39.swl.thr1_state;
thread_status[158] = `IFUPATH39.swl.thr2_state;
thread_status[159] = `IFUPATH39.swl.thr3_state;
thread_status[160] = `IFUPATH40.swl.thr0_state;
thread_status[161] = `IFUPATH40.swl.thr1_state;
thread_status[162] = `IFUPATH40.swl.thr2_state;
thread_status[163] = `IFUPATH40.swl.thr3_state;
thread_status[164] = `IFUPATH41.swl.thr0_state;
thread_status[165] = `IFUPATH41.swl.thr1_state;
thread_status[166] = `IFUPATH41.swl.thr2_state;
thread_status[167] = `IFUPATH41.swl.thr3_state;
thread_status[168] = `IFUPATH42.swl.thr0_state;
thread_status[169] = `IFUPATH42.swl.thr1_state;
thread_status[170] = `IFUPATH42.swl.thr2_state;
thread_status[171] = `IFUPATH42.swl.thr3_state;
thread_status[172] = `IFUPATH43.swl.thr0_state;
thread_status[173] = `IFUPATH43.swl.thr1_state;
thread_status[174] = `IFUPATH43.swl.thr2_state;
thread_status[175] = `IFUPATH43.swl.thr3_state;
thread_status[176] = `IFUPATH44.swl.thr0_state;
thread_status[177] = `IFUPATH44.swl.thr1_state;
thread_status[178] = `IFUPATH44.swl.thr2_state;
thread_status[179] = `IFUPATH44.swl.thr3_state;
thread_status[180] = `IFUPATH45.swl.thr0_state;
thread_status[181] = `IFUPATH45.swl.thr1_state;
thread_status[182] = `IFUPATH45.swl.thr2_state;
thread_status[183] = `IFUPATH45.swl.thr3_state;
thread_status[184] = `IFUPATH46.swl.thr0_state;
thread_status[185] = `IFUPATH46.swl.thr1_state;
thread_status[186] = `IFUPATH46.swl.thr2_state;
thread_status[187] = `IFUPATH46.swl.thr3_state;
thread_status[188] = `IFUPATH47.swl.thr0_state;
thread_status[189] = `IFUPATH47.swl.thr1_state;
thread_status[190] = `IFUPATH47.swl.thr2_state;
thread_status[191] = `IFUPATH47.swl.thr3_state;
thread_status[192] = `IFUPATH48.swl.thr0_state;
thread_status[193] = `IFUPATH48.swl.thr1_state;
thread_status[194] = `IFUPATH48.swl.thr2_state;
thread_status[195] = `IFUPATH48.swl.thr3_state;
thread_status[196] = `IFUPATH49.swl.thr0_state;
thread_status[197] = `IFUPATH49.swl.thr1_state;
thread_status[198] = `IFUPATH49.swl.thr2_state;
thread_status[199] = `IFUPATH49.swl.thr3_state;
thread_status[200] = `IFUPATH50.swl.thr0_state;
thread_status[201] = `IFUPATH50.swl.thr1_state;
thread_status[202] = `IFUPATH50.swl.thr2_state;
thread_status[203] = `IFUPATH50.swl.thr3_state;
thread_status[204] = `IFUPATH51.swl.thr0_state;
thread_status[205] = `IFUPATH51.swl.thr1_state;
thread_status[206] = `IFUPATH51.swl.thr2_state;
thread_status[207] = `IFUPATH51.swl.thr3_state;
thread_status[208] = `IFUPATH52.swl.thr0_state;
thread_status[209] = `IFUPATH52.swl.thr1_state;
thread_status[210] = `IFUPATH52.swl.thr2_state;
thread_status[211] = `IFUPATH52.swl.thr3_state;
thread_status[212] = `IFUPATH53.swl.thr0_state;
thread_status[213] = `IFUPATH53.swl.thr1_state;
thread_status[214] = `IFUPATH53.swl.thr2_state;
thread_status[215] = `IFUPATH53.swl.thr3_state;
thread_status[216] = `IFUPATH54.swl.thr0_state;
thread_status[217] = `IFUPATH54.swl.thr1_state;
thread_status[218] = `IFUPATH54.swl.thr2_state;
thread_status[219] = `IFUPATH54.swl.thr3_state;
thread_status[220] = `IFUPATH55.swl.thr0_state;
thread_status[221] = `IFUPATH55.swl.thr1_state;
thread_status[222] = `IFUPATH55.swl.thr2_state;
thread_status[223] = `IFUPATH55.swl.thr3_state;
thread_status[224] = `IFUPATH56.swl.thr0_state;
thread_status[225] = `IFUPATH56.swl.thr1_state;
thread_status[226] = `IFUPATH56.swl.thr2_state;
thread_status[227] = `IFUPATH56.swl.thr3_state;
thread_status[228] = `IFUPATH57.swl.thr0_state;
thread_status[229] = `IFUPATH57.swl.thr1_state;
thread_status[230] = `IFUPATH57.swl.thr2_state;
thread_status[231] = `IFUPATH57.swl.thr3_state;
thread_status[232] = `IFUPATH58.swl.thr0_state;
thread_status[233] = `IFUPATH58.swl.thr1_state;
thread_status[234] = `IFUPATH58.swl.thr2_state;
thread_status[235] = `IFUPATH58.swl.thr3_state;
thread_status[236] = `IFUPATH59.swl.thr0_state;
thread_status[237] = `IFUPATH59.swl.thr1_state;
thread_status[238] = `IFUPATH59.swl.thr2_state;
thread_status[239] = `IFUPATH59.swl.thr3_state;
thread_status[240] = `IFUPATH60.swl.thr0_state;
thread_status[241] = `IFUPATH60.swl.thr1_state;
thread_status[242] = `IFUPATH60.swl.thr2_state;
thread_status[243] = `IFUPATH60.swl.thr3_state;
thread_status[244] = `IFUPATH61.swl.thr0_state;
thread_status[245] = `IFUPATH61.swl.thr1_state;
thread_status[246] = `IFUPATH61.swl.thr2_state;
thread_status[247] = `IFUPATH61.swl.thr3_state;
thread_status[248] = `IFUPATH62.swl.thr0_state;
thread_status[249] = `IFUPATH62.swl.thr1_state;
thread_status[250] = `IFUPATH62.swl.thr2_state;
thread_status[251] = `IFUPATH62.swl.thr3_state;
thread_status[252] = `IFUPATH63.swl.thr0_state;
thread_status[253] = `IFUPATH63.swl.thr1_state;
thread_status[254] = `IFUPATH63.swl.thr2_state;
thread_status[255] = `IFUPATH63.swl.thr3_state;
thread_status[256] = `IFUPATH64.swl.thr0_state;
thread_status[257] = `IFUPATH64.swl.thr1_state;
thread_status[258] = `IFUPATH64.swl.thr2_state;
thread_status[259] = `IFUPATH64.swl.thr3_state;
thread_status[260] = `IFUPATH65.swl.thr0_state;
thread_status[261] = `IFUPATH65.swl.thr1_state;
thread_status[262] = `IFUPATH65.swl.thr2_state;
thread_status[263] = `IFUPATH65.swl.thr3_state;
thread_status[264] = `IFUPATH66.swl.thr0_state;
thread_status[265] = `IFUPATH66.swl.thr1_state;
thread_status[266] = `IFUPATH66.swl.thr2_state;
thread_status[267] = `IFUPATH66.swl.thr3_state;
thread_status[268] = `IFUPATH67.swl.thr0_state;
thread_status[269] = `IFUPATH67.swl.thr1_state;
thread_status[270] = `IFUPATH67.swl.thr2_state;
thread_status[271] = `IFUPATH67.swl.thr3_state;
thread_status[272] = `IFUPATH68.swl.thr0_state;
thread_status[273] = `IFUPATH68.swl.thr1_state;
thread_status[274] = `IFUPATH68.swl.thr2_state;
thread_status[275] = `IFUPATH68.swl.thr3_state;
thread_status[276] = `IFUPATH69.swl.thr0_state;
thread_status[277] = `IFUPATH69.swl.thr1_state;
thread_status[278] = `IFUPATH69.swl.thr2_state;
thread_status[279] = `IFUPATH69.swl.thr3_state;
thread_status[280] = `IFUPATH70.swl.thr0_state;
thread_status[281] = `IFUPATH70.swl.thr1_state;
thread_status[282] = `IFUPATH70.swl.thr2_state;
thread_status[283] = `IFUPATH70.swl.thr3_state;
thread_status[284] = `IFUPATH71.swl.thr0_state;
thread_status[285] = `IFUPATH71.swl.thr1_state;
thread_status[286] = `IFUPATH71.swl.thr2_state;
thread_status[287] = `IFUPATH71.swl.thr3_state;
thread_status[288] = `IFUPATH72.swl.thr0_state;
thread_status[289] = `IFUPATH72.swl.thr1_state;
thread_status[290] = `IFUPATH72.swl.thr2_state;
thread_status[291] = `IFUPATH72.swl.thr3_state;
thread_status[292] = `IFUPATH73.swl.thr0_state;
thread_status[293] = `IFUPATH73.swl.thr1_state;
thread_status[294] = `IFUPATH73.swl.thr2_state;
thread_status[295] = `IFUPATH73.swl.thr3_state;
thread_status[296] = `IFUPATH74.swl.thr0_state;
thread_status[297] = `IFUPATH74.swl.thr1_state;
thread_status[298] = `IFUPATH74.swl.thr2_state;
thread_status[299] = `IFUPATH74.swl.thr3_state;
thread_status[300] = `IFUPATH75.swl.thr0_state;
thread_status[301] = `IFUPATH75.swl.thr1_state;
thread_status[302] = `IFUPATH75.swl.thr2_state;
thread_status[303] = `IFUPATH75.swl.thr3_state;
thread_status[304] = `IFUPATH76.swl.thr0_state;
thread_status[305] = `IFUPATH76.swl.thr1_state;
thread_status[306] = `IFUPATH76.swl.thr2_state;
thread_status[307] = `IFUPATH76.swl.thr3_state;
thread_status[308] = `IFUPATH77.swl.thr0_state;
thread_status[309] = `IFUPATH77.swl.thr1_state;
thread_status[310] = `IFUPATH77.swl.thr2_state;
thread_status[311] = `IFUPATH77.swl.thr3_state;
thread_status[312] = `IFUPATH78.swl.thr0_state;
thread_status[313] = `IFUPATH78.swl.thr1_state;
thread_status[314] = `IFUPATH78.swl.thr2_state;
thread_status[315] = `IFUPATH78.swl.thr3_state;
thread_status[316] = `IFUPATH79.swl.thr0_state;
thread_status[317] = `IFUPATH79.swl.thr1_state;
thread_status[318] = `IFUPATH79.swl.thr2_state;
thread_status[319] = `IFUPATH79.swl.thr3_state;
thread_status[320] = `IFUPATH80.swl.thr0_state;
thread_status[321] = `IFUPATH80.swl.thr1_state;
thread_status[322] = `IFUPATH80.swl.thr2_state;
thread_status[323] = `IFUPATH80.swl.thr3_state;
thread_status[324] = `IFUPATH81.swl.thr0_state;
thread_status[325] = `IFUPATH81.swl.thr1_state;
thread_status[326] = `IFUPATH81.swl.thr2_state;
thread_status[327] = `IFUPATH81.swl.thr3_state;
thread_status[328] = `IFUPATH82.swl.thr0_state;
thread_status[329] = `IFUPATH82.swl.thr1_state;
thread_status[330] = `IFUPATH82.swl.thr2_state;
thread_status[331] = `IFUPATH82.swl.thr3_state;
thread_status[332] = `IFUPATH83.swl.thr0_state;
thread_status[333] = `IFUPATH83.swl.thr1_state;
thread_status[334] = `IFUPATH83.swl.thr2_state;
thread_status[335] = `IFUPATH83.swl.thr3_state;
thread_status[336] = `IFUPATH84.swl.thr0_state;
thread_status[337] = `IFUPATH84.swl.thr1_state;
thread_status[338] = `IFUPATH84.swl.thr2_state;
thread_status[339] = `IFUPATH84.swl.thr3_state;
thread_status[340] = `IFUPATH85.swl.thr0_state;
thread_status[341] = `IFUPATH85.swl.thr1_state;
thread_status[342] = `IFUPATH85.swl.thr2_state;
thread_status[343] = `IFUPATH85.swl.thr3_state;
thread_status[344] = `IFUPATH86.swl.thr0_state;
thread_status[345] = `IFUPATH86.swl.thr1_state;
thread_status[346] = `IFUPATH86.swl.thr2_state;
thread_status[347] = `IFUPATH86.swl.thr3_state;
thread_status[348] = `IFUPATH87.swl.thr0_state;
thread_status[349] = `IFUPATH87.swl.thr1_state;
thread_status[350] = `IFUPATH87.swl.thr2_state;
thread_status[351] = `IFUPATH87.swl.thr3_state;
thread_status[352] = `IFUPATH88.swl.thr0_state;
thread_status[353] = `IFUPATH88.swl.thr1_state;
thread_status[354] = `IFUPATH88.swl.thr2_state;
thread_status[355] = `IFUPATH88.swl.thr3_state;
thread_status[356] = `IFUPATH89.swl.thr0_state;
thread_status[357] = `IFUPATH89.swl.thr1_state;
thread_status[358] = `IFUPATH89.swl.thr2_state;
thread_status[359] = `IFUPATH89.swl.thr3_state;
thread_status[360] = `IFUPATH90.swl.thr0_state;
thread_status[361] = `IFUPATH90.swl.thr1_state;
thread_status[362] = `IFUPATH90.swl.thr2_state;
thread_status[363] = `IFUPATH90.swl.thr3_state;
thread_status[364] = `IFUPATH91.swl.thr0_state;
thread_status[365] = `IFUPATH91.swl.thr1_state;
thread_status[366] = `IFUPATH91.swl.thr2_state;
thread_status[367] = `IFUPATH91.swl.thr3_state;
thread_status[368] = `IFUPATH92.swl.thr0_state;
thread_status[369] = `IFUPATH92.swl.thr1_state;
thread_status[370] = `IFUPATH92.swl.thr2_state;
thread_status[371] = `IFUPATH92.swl.thr3_state;
thread_status[372] = `IFUPATH93.swl.thr0_state;
thread_status[373] = `IFUPATH93.swl.thr1_state;
thread_status[374] = `IFUPATH93.swl.thr2_state;
thread_status[375] = `IFUPATH93.swl.thr3_state;
thread_status[376] = `IFUPATH94.swl.thr0_state;
thread_status[377] = `IFUPATH94.swl.thr1_state;
thread_status[378] = `IFUPATH94.swl.thr2_state;
thread_status[379] = `IFUPATH94.swl.thr3_state;
thread_status[380] = `IFUPATH95.swl.thr0_state;
thread_status[381] = `IFUPATH95.swl.thr1_state;
thread_status[382] = `IFUPATH95.swl.thr2_state;
thread_status[383] = `IFUPATH95.swl.thr3_state;
thread_status[384] = `IFUPATH96.swl.thr0_state;
thread_status[385] = `IFUPATH96.swl.thr1_state;
thread_status[386] = `IFUPATH96.swl.thr2_state;
thread_status[387] = `IFUPATH96.swl.thr3_state;
thread_status[388] = `IFUPATH97.swl.thr0_state;
thread_status[389] = `IFUPATH97.swl.thr1_state;
thread_status[390] = `IFUPATH97.swl.thr2_state;
thread_status[391] = `IFUPATH97.swl.thr3_state;
thread_status[392] = `IFUPATH98.swl.thr0_state;
thread_status[393] = `IFUPATH98.swl.thr1_state;
thread_status[394] = `IFUPATH98.swl.thr2_state;
thread_status[395] = `IFUPATH98.swl.thr3_state;
thread_status[396] = `IFUPATH99.swl.thr0_state;
thread_status[397] = `IFUPATH99.swl.thr1_state;
thread_status[398] = `IFUPATH99.swl.thr2_state;
thread_status[399] = `IFUPATH99.swl.thr3_state;
thread_status[400] = `IFUPATH100.swl.thr0_state;
thread_status[401] = `IFUPATH100.swl.thr1_state;
thread_status[402] = `IFUPATH100.swl.thr2_state;
thread_status[403] = `IFUPATH100.swl.thr3_state;
thread_status[404] = `IFUPATH101.swl.thr0_state;
thread_status[405] = `IFUPATH101.swl.thr1_state;
thread_status[406] = `IFUPATH101.swl.thr2_state;
thread_status[407] = `IFUPATH101.swl.thr3_state;
thread_status[408] = `IFUPATH102.swl.thr0_state;
thread_status[409] = `IFUPATH102.swl.thr1_state;
thread_status[410] = `IFUPATH102.swl.thr2_state;
thread_status[411] = `IFUPATH102.swl.thr3_state;
thread_status[412] = `IFUPATH103.swl.thr0_state;
thread_status[413] = `IFUPATH103.swl.thr1_state;
thread_status[414] = `IFUPATH103.swl.thr2_state;
thread_status[415] = `IFUPATH103.swl.thr3_state;
thread_status[416] = `IFUPATH104.swl.thr0_state;
thread_status[417] = `IFUPATH104.swl.thr1_state;
thread_status[418] = `IFUPATH104.swl.thr2_state;
thread_status[419] = `IFUPATH104.swl.thr3_state;
thread_status[420] = `IFUPATH105.swl.thr0_state;
thread_status[421] = `IFUPATH105.swl.thr1_state;
thread_status[422] = `IFUPATH105.swl.thr2_state;
thread_status[423] = `IFUPATH105.swl.thr3_state;
thread_status[424] = `IFUPATH106.swl.thr0_state;
thread_status[425] = `IFUPATH106.swl.thr1_state;
thread_status[426] = `IFUPATH106.swl.thr2_state;
thread_status[427] = `IFUPATH106.swl.thr3_state;
thread_status[428] = `IFUPATH107.swl.thr0_state;
thread_status[429] = `IFUPATH107.swl.thr1_state;
thread_status[430] = `IFUPATH107.swl.thr2_state;
thread_status[431] = `IFUPATH107.swl.thr3_state;
thread_status[432] = `IFUPATH108.swl.thr0_state;
thread_status[433] = `IFUPATH108.swl.thr1_state;
thread_status[434] = `IFUPATH108.swl.thr2_state;
thread_status[435] = `IFUPATH108.swl.thr3_state;
thread_status[436] = `IFUPATH109.swl.thr0_state;
thread_status[437] = `IFUPATH109.swl.thr1_state;
thread_status[438] = `IFUPATH109.swl.thr2_state;
thread_status[439] = `IFUPATH109.swl.thr3_state;
thread_status[440] = `IFUPATH110.swl.thr0_state;
thread_status[441] = `IFUPATH110.swl.thr1_state;
thread_status[442] = `IFUPATH110.swl.thr2_state;
thread_status[443] = `IFUPATH110.swl.thr3_state;
thread_status[444] = `IFUPATH111.swl.thr0_state;
thread_status[445] = `IFUPATH111.swl.thr1_state;
thread_status[446] = `IFUPATH111.swl.thr2_state;
thread_status[447] = `IFUPATH111.swl.thr3_state;
thread_status[448] = `IFUPATH112.swl.thr0_state;
thread_status[449] = `IFUPATH112.swl.thr1_state;
thread_status[450] = `IFUPATH112.swl.thr2_state;
thread_status[451] = `IFUPATH112.swl.thr3_state;
thread_status[452] = `IFUPATH113.swl.thr0_state;
thread_status[453] = `IFUPATH113.swl.thr1_state;
thread_status[454] = `IFUPATH113.swl.thr2_state;
thread_status[455] = `IFUPATH113.swl.thr3_state;
thread_status[456] = `IFUPATH114.swl.thr0_state;
thread_status[457] = `IFUPATH114.swl.thr1_state;
thread_status[458] = `IFUPATH114.swl.thr2_state;
thread_status[459] = `IFUPATH114.swl.thr3_state;
thread_status[460] = `IFUPATH115.swl.thr0_state;
thread_status[461] = `IFUPATH115.swl.thr1_state;
thread_status[462] = `IFUPATH115.swl.thr2_state;
thread_status[463] = `IFUPATH115.swl.thr3_state;
thread_status[464] = `IFUPATH116.swl.thr0_state;
thread_status[465] = `IFUPATH116.swl.thr1_state;
thread_status[466] = `IFUPATH116.swl.thr2_state;
thread_status[467] = `IFUPATH116.swl.thr3_state;
thread_status[468] = `IFUPATH117.swl.thr0_state;
thread_status[469] = `IFUPATH117.swl.thr1_state;
thread_status[470] = `IFUPATH117.swl.thr2_state;
thread_status[471] = `IFUPATH117.swl.thr3_state;
thread_status[472] = `IFUPATH118.swl.thr0_state;
thread_status[473] = `IFUPATH118.swl.thr1_state;
thread_status[474] = `IFUPATH118.swl.thr2_state;
thread_status[475] = `IFUPATH118.swl.thr3_state;
thread_status[476] = `IFUPATH119.swl.thr0_state;
thread_status[477] = `IFUPATH119.swl.thr1_state;
thread_status[478] = `IFUPATH119.swl.thr2_state;
thread_status[479] = `IFUPATH119.swl.thr3_state;
thread_status[480] = `IFUPATH120.swl.thr0_state;
thread_status[481] = `IFUPATH120.swl.thr1_state;
thread_status[482] = `IFUPATH120.swl.thr2_state;
thread_status[483] = `IFUPATH120.swl.thr3_state;
thread_status[484] = `IFUPATH121.swl.thr0_state;
thread_status[485] = `IFUPATH121.swl.thr1_state;
thread_status[486] = `IFUPATH121.swl.thr2_state;
thread_status[487] = `IFUPATH121.swl.thr3_state;
thread_status[488] = `IFUPATH122.swl.thr0_state;
thread_status[489] = `IFUPATH122.swl.thr1_state;
thread_status[490] = `IFUPATH122.swl.thr2_state;
thread_status[491] = `IFUPATH122.swl.thr3_state;
thread_status[492] = `IFUPATH123.swl.thr0_state;
thread_status[493] = `IFUPATH123.swl.thr1_state;
thread_status[494] = `IFUPATH123.swl.thr2_state;
thread_status[495] = `IFUPATH123.swl.thr3_state;
thread_status[496] = `IFUPATH124.swl.thr0_state;
thread_status[497] = `IFUPATH124.swl.thr1_state;
thread_status[498] = `IFUPATH124.swl.thr2_state;
thread_status[499] = `IFUPATH124.swl.thr3_state;
thread_status[500] = `IFUPATH125.swl.thr0_state;
thread_status[501] = `IFUPATH125.swl.thr1_state;
thread_status[502] = `IFUPATH125.swl.thr2_state;
thread_status[503] = `IFUPATH125.swl.thr3_state;
thread_status[504] = `IFUPATH126.swl.thr0_state;
thread_status[505] = `IFUPATH126.swl.thr1_state;
thread_status[506] = `IFUPATH126.swl.thr2_state;
thread_status[507] = `IFUPATH126.swl.thr3_state;
thread_status[508] = `IFUPATH127.swl.thr0_state;
thread_status[509] = `IFUPATH127.swl.thr1_state;
thread_status[510] = `IFUPATH127.swl.thr2_state;
thread_status[511] = `IFUPATH127.swl.thr3_state;
thread_status[512] = `IFUPATH128.swl.thr0_state;
thread_status[513] = `IFUPATH128.swl.thr1_state;
thread_status[514] = `IFUPATH128.swl.thr2_state;
thread_status[515] = `IFUPATH128.swl.thr3_state;
thread_status[516] = `IFUPATH129.swl.thr0_state;
thread_status[517] = `IFUPATH129.swl.thr1_state;
thread_status[518] = `IFUPATH129.swl.thr2_state;
thread_status[519] = `IFUPATH129.swl.thr3_state;
thread_status[520] = `IFUPATH130.swl.thr0_state;
thread_status[521] = `IFUPATH130.swl.thr1_state;
thread_status[522] = `IFUPATH130.swl.thr2_state;
thread_status[523] = `IFUPATH130.swl.thr3_state;
thread_status[524] = `IFUPATH131.swl.thr0_state;
thread_status[525] = `IFUPATH131.swl.thr1_state;
thread_status[526] = `IFUPATH131.swl.thr2_state;
thread_status[527] = `IFUPATH131.swl.thr3_state;
thread_status[528] = `IFUPATH132.swl.thr0_state;
thread_status[529] = `IFUPATH132.swl.thr1_state;
thread_status[530] = `IFUPATH132.swl.thr2_state;
thread_status[531] = `IFUPATH132.swl.thr3_state;
thread_status[532] = `IFUPATH133.swl.thr0_state;
thread_status[533] = `IFUPATH133.swl.thr1_state;
thread_status[534] = `IFUPATH133.swl.thr2_state;
thread_status[535] = `IFUPATH133.swl.thr3_state;
thread_status[536] = `IFUPATH134.swl.thr0_state;
thread_status[537] = `IFUPATH134.swl.thr1_state;
thread_status[538] = `IFUPATH134.swl.thr2_state;
thread_status[539] = `IFUPATH134.swl.thr3_state;
thread_status[540] = `IFUPATH135.swl.thr0_state;
thread_status[541] = `IFUPATH135.swl.thr1_state;
thread_status[542] = `IFUPATH135.swl.thr2_state;
thread_status[543] = `IFUPATH135.swl.thr3_state;
thread_status[544] = `IFUPATH136.swl.thr0_state;
thread_status[545] = `IFUPATH136.swl.thr1_state;
thread_status[546] = `IFUPATH136.swl.thr2_state;
thread_status[547] = `IFUPATH136.swl.thr3_state;
thread_status[548] = `IFUPATH137.swl.thr0_state;
thread_status[549] = `IFUPATH137.swl.thr1_state;
thread_status[550] = `IFUPATH137.swl.thr2_state;
thread_status[551] = `IFUPATH137.swl.thr3_state;
thread_status[552] = `IFUPATH138.swl.thr0_state;
thread_status[553] = `IFUPATH138.swl.thr1_state;
thread_status[554] = `IFUPATH138.swl.thr2_state;
thread_status[555] = `IFUPATH138.swl.thr3_state;
thread_status[556] = `IFUPATH139.swl.thr0_state;
thread_status[557] = `IFUPATH139.swl.thr1_state;
thread_status[558] = `IFUPATH139.swl.thr2_state;
thread_status[559] = `IFUPATH139.swl.thr3_state;
thread_status[560] = `IFUPATH140.swl.thr0_state;
thread_status[561] = `IFUPATH140.swl.thr1_state;
thread_status[562] = `IFUPATH140.swl.thr2_state;
thread_status[563] = `IFUPATH140.swl.thr3_state;
thread_status[564] = `IFUPATH141.swl.thr0_state;
thread_status[565] = `IFUPATH141.swl.thr1_state;
thread_status[566] = `IFUPATH141.swl.thr2_state;
thread_status[567] = `IFUPATH141.swl.thr3_state;
thread_status[568] = `IFUPATH142.swl.thr0_state;
thread_status[569] = `IFUPATH142.swl.thr1_state;
thread_status[570] = `IFUPATH142.swl.thr2_state;
thread_status[571] = `IFUPATH142.swl.thr3_state;
thread_status[572] = `IFUPATH143.swl.thr0_state;
thread_status[573] = `IFUPATH143.swl.thr1_state;
thread_status[574] = `IFUPATH143.swl.thr2_state;
thread_status[575] = `IFUPATH143.swl.thr3_state;
thread_status[576] = `IFUPATH144.swl.thr0_state;
thread_status[577] = `IFUPATH144.swl.thr1_state;
thread_status[578] = `IFUPATH144.swl.thr2_state;
thread_status[579] = `IFUPATH144.swl.thr3_state;
thread_status[580] = `IFUPATH145.swl.thr0_state;
thread_status[581] = `IFUPATH145.swl.thr1_state;
thread_status[582] = `IFUPATH145.swl.thr2_state;
thread_status[583] = `IFUPATH145.swl.thr3_state;
thread_status[584] = `IFUPATH146.swl.thr0_state;
thread_status[585] = `IFUPATH146.swl.thr1_state;
thread_status[586] = `IFUPATH146.swl.thr2_state;
thread_status[587] = `IFUPATH146.swl.thr3_state;
thread_status[588] = `IFUPATH147.swl.thr0_state;
thread_status[589] = `IFUPATH147.swl.thr1_state;
thread_status[590] = `IFUPATH147.swl.thr2_state;
thread_status[591] = `IFUPATH147.swl.thr3_state;
thread_status[592] = `IFUPATH148.swl.thr0_state;
thread_status[593] = `IFUPATH148.swl.thr1_state;
thread_status[594] = `IFUPATH148.swl.thr2_state;
thread_status[595] = `IFUPATH148.swl.thr3_state;
thread_status[596] = `IFUPATH149.swl.thr0_state;
thread_status[597] = `IFUPATH149.swl.thr1_state;
thread_status[598] = `IFUPATH149.swl.thr2_state;
thread_status[599] = `IFUPATH149.swl.thr3_state;
thread_status[600] = `IFUPATH150.swl.thr0_state;
thread_status[601] = `IFUPATH150.swl.thr1_state;
thread_status[602] = `IFUPATH150.swl.thr2_state;
thread_status[603] = `IFUPATH150.swl.thr3_state;
thread_status[604] = `IFUPATH151.swl.thr0_state;
thread_status[605] = `IFUPATH151.swl.thr1_state;
thread_status[606] = `IFUPATH151.swl.thr2_state;
thread_status[607] = `IFUPATH151.swl.thr3_state;
thread_status[608] = `IFUPATH152.swl.thr0_state;
thread_status[609] = `IFUPATH152.swl.thr1_state;
thread_status[610] = `IFUPATH152.swl.thr2_state;
thread_status[611] = `IFUPATH152.swl.thr3_state;
thread_status[612] = `IFUPATH153.swl.thr0_state;
thread_status[613] = `IFUPATH153.swl.thr1_state;
thread_status[614] = `IFUPATH153.swl.thr2_state;
thread_status[615] = `IFUPATH153.swl.thr3_state;
thread_status[616] = `IFUPATH154.swl.thr0_state;
thread_status[617] = `IFUPATH154.swl.thr1_state;
thread_status[618] = `IFUPATH154.swl.thr2_state;
thread_status[619] = `IFUPATH154.swl.thr3_state;
thread_status[620] = `IFUPATH155.swl.thr0_state;
thread_status[621] = `IFUPATH155.swl.thr1_state;
thread_status[622] = `IFUPATH155.swl.thr2_state;
thread_status[623] = `IFUPATH155.swl.thr3_state;
thread_status[624] = `IFUPATH156.swl.thr0_state;
thread_status[625] = `IFUPATH156.swl.thr1_state;
thread_status[626] = `IFUPATH156.swl.thr2_state;
thread_status[627] = `IFUPATH156.swl.thr3_state;
thread_status[628] = `IFUPATH157.swl.thr0_state;
thread_status[629] = `IFUPATH157.swl.thr1_state;
thread_status[630] = `IFUPATH157.swl.thr2_state;
thread_status[631] = `IFUPATH157.swl.thr3_state;
thread_status[632] = `IFUPATH158.swl.thr0_state;
thread_status[633] = `IFUPATH158.swl.thr1_state;
thread_status[634] = `IFUPATH158.swl.thr2_state;
thread_status[635] = `IFUPATH158.swl.thr3_state;
thread_status[636] = `IFUPATH159.swl.thr0_state;
thread_status[637] = `IFUPATH159.swl.thr1_state;
thread_status[638] = `IFUPATH159.swl.thr2_state;
thread_status[639] = `IFUPATH159.swl.thr3_state;
thread_status[640] = `IFUPATH160.swl.thr0_state;
thread_status[641] = `IFUPATH160.swl.thr1_state;
thread_status[642] = `IFUPATH160.swl.thr2_state;
thread_status[643] = `IFUPATH160.swl.thr3_state;
thread_status[644] = `IFUPATH161.swl.thr0_state;
thread_status[645] = `IFUPATH161.swl.thr1_state;
thread_status[646] = `IFUPATH161.swl.thr2_state;
thread_status[647] = `IFUPATH161.swl.thr3_state;
thread_status[648] = `IFUPATH162.swl.thr0_state;
thread_status[649] = `IFUPATH162.swl.thr1_state;
thread_status[650] = `IFUPATH162.swl.thr2_state;
thread_status[651] = `IFUPATH162.swl.thr3_state;
thread_status[652] = `IFUPATH163.swl.thr0_state;
thread_status[653] = `IFUPATH163.swl.thr1_state;
thread_status[654] = `IFUPATH163.swl.thr2_state;
thread_status[655] = `IFUPATH163.swl.thr3_state;
thread_status[656] = `IFUPATH164.swl.thr0_state;
thread_status[657] = `IFUPATH164.swl.thr1_state;
thread_status[658] = `IFUPATH164.swl.thr2_state;
thread_status[659] = `IFUPATH164.swl.thr3_state;
thread_status[660] = `IFUPATH165.swl.thr0_state;
thread_status[661] = `IFUPATH165.swl.thr1_state;
thread_status[662] = `IFUPATH165.swl.thr2_state;
thread_status[663] = `IFUPATH165.swl.thr3_state;
thread_status[664] = `IFUPATH166.swl.thr0_state;
thread_status[665] = `IFUPATH166.swl.thr1_state;
thread_status[666] = `IFUPATH166.swl.thr2_state;
thread_status[667] = `IFUPATH166.swl.thr3_state;
thread_status[668] = `IFUPATH167.swl.thr0_state;
thread_status[669] = `IFUPATH167.swl.thr1_state;
thread_status[670] = `IFUPATH167.swl.thr2_state;
thread_status[671] = `IFUPATH167.swl.thr3_state;
thread_status[672] = `IFUPATH168.swl.thr0_state;
thread_status[673] = `IFUPATH168.swl.thr1_state;
thread_status[674] = `IFUPATH168.swl.thr2_state;
thread_status[675] = `IFUPATH168.swl.thr3_state;
thread_status[676] = `IFUPATH169.swl.thr0_state;
thread_status[677] = `IFUPATH169.swl.thr1_state;
thread_status[678] = `IFUPATH169.swl.thr2_state;
thread_status[679] = `IFUPATH169.swl.thr3_state;
thread_status[680] = `IFUPATH170.swl.thr0_state;
thread_status[681] = `IFUPATH170.swl.thr1_state;
thread_status[682] = `IFUPATH170.swl.thr2_state;
thread_status[683] = `IFUPATH170.swl.thr3_state;
thread_status[684] = `IFUPATH171.swl.thr0_state;
thread_status[685] = `IFUPATH171.swl.thr1_state;
thread_status[686] = `IFUPATH171.swl.thr2_state;
thread_status[687] = `IFUPATH171.swl.thr3_state;
thread_status[688] = `IFUPATH172.swl.thr0_state;
thread_status[689] = `IFUPATH172.swl.thr1_state;
thread_status[690] = `IFUPATH172.swl.thr2_state;
thread_status[691] = `IFUPATH172.swl.thr3_state;
thread_status[692] = `IFUPATH173.swl.thr0_state;
thread_status[693] = `IFUPATH173.swl.thr1_state;
thread_status[694] = `IFUPATH173.swl.thr2_state;
thread_status[695] = `IFUPATH173.swl.thr3_state;
thread_status[696] = `IFUPATH174.swl.thr0_state;
thread_status[697] = `IFUPATH174.swl.thr1_state;
thread_status[698] = `IFUPATH174.swl.thr2_state;
thread_status[699] = `IFUPATH174.swl.thr3_state;
thread_status[700] = `IFUPATH175.swl.thr0_state;
thread_status[701] = `IFUPATH175.swl.thr1_state;
thread_status[702] = `IFUPATH175.swl.thr2_state;
thread_status[703] = `IFUPATH175.swl.thr3_state;
thread_status[704] = `IFUPATH176.swl.thr0_state;
thread_status[705] = `IFUPATH176.swl.thr1_state;
thread_status[706] = `IFUPATH176.swl.thr2_state;
thread_status[707] = `IFUPATH176.swl.thr3_state;
thread_status[708] = `IFUPATH177.swl.thr0_state;
thread_status[709] = `IFUPATH177.swl.thr1_state;
thread_status[710] = `IFUPATH177.swl.thr2_state;
thread_status[711] = `IFUPATH177.swl.thr3_state;
thread_status[712] = `IFUPATH178.swl.thr0_state;
thread_status[713] = `IFUPATH178.swl.thr1_state;
thread_status[714] = `IFUPATH178.swl.thr2_state;
thread_status[715] = `IFUPATH178.swl.thr3_state;
thread_status[716] = `IFUPATH179.swl.thr0_state;
thread_status[717] = `IFUPATH179.swl.thr1_state;
thread_status[718] = `IFUPATH179.swl.thr2_state;
thread_status[719] = `IFUPATH179.swl.thr3_state;
thread_status[720] = `IFUPATH180.swl.thr0_state;
thread_status[721] = `IFUPATH180.swl.thr1_state;
thread_status[722] = `IFUPATH180.swl.thr2_state;
thread_status[723] = `IFUPATH180.swl.thr3_state;
thread_status[724] = `IFUPATH181.swl.thr0_state;
thread_status[725] = `IFUPATH181.swl.thr1_state;
thread_status[726] = `IFUPATH181.swl.thr2_state;
thread_status[727] = `IFUPATH181.swl.thr3_state;
thread_status[728] = `IFUPATH182.swl.thr0_state;
thread_status[729] = `IFUPATH182.swl.thr1_state;
thread_status[730] = `IFUPATH182.swl.thr2_state;
thread_status[731] = `IFUPATH182.swl.thr3_state;
thread_status[732] = `IFUPATH183.swl.thr0_state;
thread_status[733] = `IFUPATH183.swl.thr1_state;
thread_status[734] = `IFUPATH183.swl.thr2_state;
thread_status[735] = `IFUPATH183.swl.thr3_state;
thread_status[736] = `IFUPATH184.swl.thr0_state;
thread_status[737] = `IFUPATH184.swl.thr1_state;
thread_status[738] = `IFUPATH184.swl.thr2_state;
thread_status[739] = `IFUPATH184.swl.thr3_state;
thread_status[740] = `IFUPATH185.swl.thr0_state;
thread_status[741] = `IFUPATH185.swl.thr1_state;
thread_status[742] = `IFUPATH185.swl.thr2_state;
thread_status[743] = `IFUPATH185.swl.thr3_state;
thread_status[744] = `IFUPATH186.swl.thr0_state;
thread_status[745] = `IFUPATH186.swl.thr1_state;
thread_status[746] = `IFUPATH186.swl.thr2_state;
thread_status[747] = `IFUPATH186.swl.thr3_state;
thread_status[748] = `IFUPATH187.swl.thr0_state;
thread_status[749] = `IFUPATH187.swl.thr1_state;
thread_status[750] = `IFUPATH187.swl.thr2_state;
thread_status[751] = `IFUPATH187.swl.thr3_state;
thread_status[752] = `IFUPATH188.swl.thr0_state;
thread_status[753] = `IFUPATH188.swl.thr1_state;
thread_status[754] = `IFUPATH188.swl.thr2_state;
thread_status[755] = `IFUPATH188.swl.thr3_state;
thread_status[756] = `IFUPATH189.swl.thr0_state;
thread_status[757] = `IFUPATH189.swl.thr1_state;
thread_status[758] = `IFUPATH189.swl.thr2_state;
thread_status[759] = `IFUPATH189.swl.thr3_state;
thread_status[760] = `IFUPATH190.swl.thr0_state;
thread_status[761] = `IFUPATH190.swl.thr1_state;
thread_status[762] = `IFUPATH190.swl.thr2_state;
thread_status[763] = `IFUPATH190.swl.thr3_state;
thread_status[764] = `IFUPATH191.swl.thr0_state;
thread_status[765] = `IFUPATH191.swl.thr1_state;
thread_status[766] = `IFUPATH191.swl.thr2_state;
thread_status[767] = `IFUPATH191.swl.thr3_state;
thread_status[768] = `IFUPATH192.swl.thr0_state;
thread_status[769] = `IFUPATH192.swl.thr1_state;
thread_status[770] = `IFUPATH192.swl.thr2_state;
thread_status[771] = `IFUPATH192.swl.thr3_state;
thread_status[772] = `IFUPATH193.swl.thr0_state;
thread_status[773] = `IFUPATH193.swl.thr1_state;
thread_status[774] = `IFUPATH193.swl.thr2_state;
thread_status[775] = `IFUPATH193.swl.thr3_state;
thread_status[776] = `IFUPATH194.swl.thr0_state;
thread_status[777] = `IFUPATH194.swl.thr1_state;
thread_status[778] = `IFUPATH194.swl.thr2_state;
thread_status[779] = `IFUPATH194.swl.thr3_state;
thread_status[780] = `IFUPATH195.swl.thr0_state;
thread_status[781] = `IFUPATH195.swl.thr1_state;
thread_status[782] = `IFUPATH195.swl.thr2_state;
thread_status[783] = `IFUPATH195.swl.thr3_state;
thread_status[784] = `IFUPATH196.swl.thr0_state;
thread_status[785] = `IFUPATH196.swl.thr1_state;
thread_status[786] = `IFUPATH196.swl.thr2_state;
thread_status[787] = `IFUPATH196.swl.thr3_state;
thread_status[788] = `IFUPATH197.swl.thr0_state;
thread_status[789] = `IFUPATH197.swl.thr1_state;
thread_status[790] = `IFUPATH197.swl.thr2_state;
thread_status[791] = `IFUPATH197.swl.thr3_state;
thread_status[792] = `IFUPATH198.swl.thr0_state;
thread_status[793] = `IFUPATH198.swl.thr1_state;
thread_status[794] = `IFUPATH198.swl.thr2_state;
thread_status[795] = `IFUPATH198.swl.thr3_state;
thread_status[796] = `IFUPATH199.swl.thr0_state;
thread_status[797] = `IFUPATH199.swl.thr1_state;
thread_status[798] = `IFUPATH199.swl.thr2_state;
thread_status[799] = `IFUPATH199.swl.thr3_state;
thread_status[800] = `IFUPATH200.swl.thr0_state;
thread_status[801] = `IFUPATH200.swl.thr1_state;
thread_status[802] = `IFUPATH200.swl.thr2_state;
thread_status[803] = `IFUPATH200.swl.thr3_state;
thread_status[804] = `IFUPATH201.swl.thr0_state;
thread_status[805] = `IFUPATH201.swl.thr1_state;
thread_status[806] = `IFUPATH201.swl.thr2_state;
thread_status[807] = `IFUPATH201.swl.thr3_state;
thread_status[808] = `IFUPATH202.swl.thr0_state;
thread_status[809] = `IFUPATH202.swl.thr1_state;
thread_status[810] = `IFUPATH202.swl.thr2_state;
thread_status[811] = `IFUPATH202.swl.thr3_state;
thread_status[812] = `IFUPATH203.swl.thr0_state;
thread_status[813] = `IFUPATH203.swl.thr1_state;
thread_status[814] = `IFUPATH203.swl.thr2_state;
thread_status[815] = `IFUPATH203.swl.thr3_state;
thread_status[816] = `IFUPATH204.swl.thr0_state;
thread_status[817] = `IFUPATH204.swl.thr1_state;
thread_status[818] = `IFUPATH204.swl.thr2_state;
thread_status[819] = `IFUPATH204.swl.thr3_state;
thread_status[820] = `IFUPATH205.swl.thr0_state;
thread_status[821] = `IFUPATH205.swl.thr1_state;
thread_status[822] = `IFUPATH205.swl.thr2_state;
thread_status[823] = `IFUPATH205.swl.thr3_state;
thread_status[824] = `IFUPATH206.swl.thr0_state;
thread_status[825] = `IFUPATH206.swl.thr1_state;
thread_status[826] = `IFUPATH206.swl.thr2_state;
thread_status[827] = `IFUPATH206.swl.thr3_state;
thread_status[828] = `IFUPATH207.swl.thr0_state;
thread_status[829] = `IFUPATH207.swl.thr1_state;
thread_status[830] = `IFUPATH207.swl.thr2_state;
thread_status[831] = `IFUPATH207.swl.thr3_state;
thread_status[832] = `IFUPATH208.swl.thr0_state;
thread_status[833] = `IFUPATH208.swl.thr1_state;
thread_status[834] = `IFUPATH208.swl.thr2_state;
thread_status[835] = `IFUPATH208.swl.thr3_state;
thread_status[836] = `IFUPATH209.swl.thr0_state;
thread_status[837] = `IFUPATH209.swl.thr1_state;
thread_status[838] = `IFUPATH209.swl.thr2_state;
thread_status[839] = `IFUPATH209.swl.thr3_state;
thread_status[840] = `IFUPATH210.swl.thr0_state;
thread_status[841] = `IFUPATH210.swl.thr1_state;
thread_status[842] = `IFUPATH210.swl.thr2_state;
thread_status[843] = `IFUPATH210.swl.thr3_state;
thread_status[844] = `IFUPATH211.swl.thr0_state;
thread_status[845] = `IFUPATH211.swl.thr1_state;
thread_status[846] = `IFUPATH211.swl.thr2_state;
thread_status[847] = `IFUPATH211.swl.thr3_state;
thread_status[848] = `IFUPATH212.swl.thr0_state;
thread_status[849] = `IFUPATH212.swl.thr1_state;
thread_status[850] = `IFUPATH212.swl.thr2_state;
thread_status[851] = `IFUPATH212.swl.thr3_state;
thread_status[852] = `IFUPATH213.swl.thr0_state;
thread_status[853] = `IFUPATH213.swl.thr1_state;
thread_status[854] = `IFUPATH213.swl.thr2_state;
thread_status[855] = `IFUPATH213.swl.thr3_state;
thread_status[856] = `IFUPATH214.swl.thr0_state;
thread_status[857] = `IFUPATH214.swl.thr1_state;
thread_status[858] = `IFUPATH214.swl.thr2_state;
thread_status[859] = `IFUPATH214.swl.thr3_state;
thread_status[860] = `IFUPATH215.swl.thr0_state;
thread_status[861] = `IFUPATH215.swl.thr1_state;
thread_status[862] = `IFUPATH215.swl.thr2_state;
thread_status[863] = `IFUPATH215.swl.thr3_state;
thread_status[864] = `IFUPATH216.swl.thr0_state;
thread_status[865] = `IFUPATH216.swl.thr1_state;
thread_status[866] = `IFUPATH216.swl.thr2_state;
thread_status[867] = `IFUPATH216.swl.thr3_state;
thread_status[868] = `IFUPATH217.swl.thr0_state;
thread_status[869] = `IFUPATH217.swl.thr1_state;
thread_status[870] = `IFUPATH217.swl.thr2_state;
thread_status[871] = `IFUPATH217.swl.thr3_state;
thread_status[872] = `IFUPATH218.swl.thr0_state;
thread_status[873] = `IFUPATH218.swl.thr1_state;
thread_status[874] = `IFUPATH218.swl.thr2_state;
thread_status[875] = `IFUPATH218.swl.thr3_state;
thread_status[876] = `IFUPATH219.swl.thr0_state;
thread_status[877] = `IFUPATH219.swl.thr1_state;
thread_status[878] = `IFUPATH219.swl.thr2_state;
thread_status[879] = `IFUPATH219.swl.thr3_state;
thread_status[880] = `IFUPATH220.swl.thr0_state;
thread_status[881] = `IFUPATH220.swl.thr1_state;
thread_status[882] = `IFUPATH220.swl.thr2_state;
thread_status[883] = `IFUPATH220.swl.thr3_state;
thread_status[884] = `IFUPATH221.swl.thr0_state;
thread_status[885] = `IFUPATH221.swl.thr1_state;
thread_status[886] = `IFUPATH221.swl.thr2_state;
thread_status[887] = `IFUPATH221.swl.thr3_state;
thread_status[888] = `IFUPATH222.swl.thr0_state;
thread_status[889] = `IFUPATH222.swl.thr1_state;
thread_status[890] = `IFUPATH222.swl.thr2_state;
thread_status[891] = `IFUPATH222.swl.thr3_state;
thread_status[892] = `IFUPATH223.swl.thr0_state;
thread_status[893] = `IFUPATH223.swl.thr1_state;
thread_status[894] = `IFUPATH223.swl.thr2_state;
thread_status[895] = `IFUPATH223.swl.thr3_state;
thread_status[896] = `IFUPATH224.swl.thr0_state;
thread_status[897] = `IFUPATH224.swl.thr1_state;
thread_status[898] = `IFUPATH224.swl.thr2_state;
thread_status[899] = `IFUPATH224.swl.thr3_state;
thread_status[900] = `IFUPATH225.swl.thr0_state;
thread_status[901] = `IFUPATH225.swl.thr1_state;
thread_status[902] = `IFUPATH225.swl.thr2_state;
thread_status[903] = `IFUPATH225.swl.thr3_state;
thread_status[904] = `IFUPATH226.swl.thr0_state;
thread_status[905] = `IFUPATH226.swl.thr1_state;
thread_status[906] = `IFUPATH226.swl.thr2_state;
thread_status[907] = `IFUPATH226.swl.thr3_state;
thread_status[908] = `IFUPATH227.swl.thr0_state;
thread_status[909] = `IFUPATH227.swl.thr1_state;
thread_status[910] = `IFUPATH227.swl.thr2_state;
thread_status[911] = `IFUPATH227.swl.thr3_state;
thread_status[912] = `IFUPATH228.swl.thr0_state;
thread_status[913] = `IFUPATH228.swl.thr1_state;
thread_status[914] = `IFUPATH228.swl.thr2_state;
thread_status[915] = `IFUPATH228.swl.thr3_state;
thread_status[916] = `IFUPATH229.swl.thr0_state;
thread_status[917] = `IFUPATH229.swl.thr1_state;
thread_status[918] = `IFUPATH229.swl.thr2_state;
thread_status[919] = `IFUPATH229.swl.thr3_state;
thread_status[920] = `IFUPATH230.swl.thr0_state;
thread_status[921] = `IFUPATH230.swl.thr1_state;
thread_status[922] = `IFUPATH230.swl.thr2_state;
thread_status[923] = `IFUPATH230.swl.thr3_state;
thread_status[924] = `IFUPATH231.swl.thr0_state;
thread_status[925] = `IFUPATH231.swl.thr1_state;
thread_status[926] = `IFUPATH231.swl.thr2_state;
thread_status[927] = `IFUPATH231.swl.thr3_state;
thread_status[928] = `IFUPATH232.swl.thr0_state;
thread_status[929] = `IFUPATH232.swl.thr1_state;
thread_status[930] = `IFUPATH232.swl.thr2_state;
thread_status[931] = `IFUPATH232.swl.thr3_state;
thread_status[932] = `IFUPATH233.swl.thr0_state;
thread_status[933] = `IFUPATH233.swl.thr1_state;
thread_status[934] = `IFUPATH233.swl.thr2_state;
thread_status[935] = `IFUPATH233.swl.thr3_state;
thread_status[936] = `IFUPATH234.swl.thr0_state;
thread_status[937] = `IFUPATH234.swl.thr1_state;
thread_status[938] = `IFUPATH234.swl.thr2_state;
thread_status[939] = `IFUPATH234.swl.thr3_state;
thread_status[940] = `IFUPATH235.swl.thr0_state;
thread_status[941] = `IFUPATH235.swl.thr1_state;
thread_status[942] = `IFUPATH235.swl.thr2_state;
thread_status[943] = `IFUPATH235.swl.thr3_state;
thread_status[944] = `IFUPATH236.swl.thr0_state;
thread_status[945] = `IFUPATH236.swl.thr1_state;
thread_status[946] = `IFUPATH236.swl.thr2_state;
thread_status[947] = `IFUPATH236.swl.thr3_state;
thread_status[948] = `IFUPATH237.swl.thr0_state;
thread_status[949] = `IFUPATH237.swl.thr1_state;
thread_status[950] = `IFUPATH237.swl.thr2_state;
thread_status[951] = `IFUPATH237.swl.thr3_state;
thread_status[952] = `IFUPATH238.swl.thr0_state;
thread_status[953] = `IFUPATH238.swl.thr1_state;
thread_status[954] = `IFUPATH238.swl.thr2_state;
thread_status[955] = `IFUPATH238.swl.thr3_state;
thread_status[956] = `IFUPATH239.swl.thr0_state;
thread_status[957] = `IFUPATH239.swl.thr1_state;
thread_status[958] = `IFUPATH239.swl.thr2_state;
thread_status[959] = `IFUPATH239.swl.thr3_state;
thread_status[960] = `IFUPATH240.swl.thr0_state;
thread_status[961] = `IFUPATH240.swl.thr1_state;
thread_status[962] = `IFUPATH240.swl.thr2_state;
thread_status[963] = `IFUPATH240.swl.thr3_state;
thread_status[964] = `IFUPATH241.swl.thr0_state;
thread_status[965] = `IFUPATH241.swl.thr1_state;
thread_status[966] = `IFUPATH241.swl.thr2_state;
thread_status[967] = `IFUPATH241.swl.thr3_state;
thread_status[968] = `IFUPATH242.swl.thr0_state;
thread_status[969] = `IFUPATH242.swl.thr1_state;
thread_status[970] = `IFUPATH242.swl.thr2_state;
thread_status[971] = `IFUPATH242.swl.thr3_state;
thread_status[972] = `IFUPATH243.swl.thr0_state;
thread_status[973] = `IFUPATH243.swl.thr1_state;
thread_status[974] = `IFUPATH243.swl.thr2_state;
thread_status[975] = `IFUPATH243.swl.thr3_state;
thread_status[976] = `IFUPATH244.swl.thr0_state;
thread_status[977] = `IFUPATH244.swl.thr1_state;
thread_status[978] = `IFUPATH244.swl.thr2_state;
thread_status[979] = `IFUPATH244.swl.thr3_state;
thread_status[980] = `IFUPATH245.swl.thr0_state;
thread_status[981] = `IFUPATH245.swl.thr1_state;
thread_status[982] = `IFUPATH245.swl.thr2_state;
thread_status[983] = `IFUPATH245.swl.thr3_state;
thread_status[984] = `IFUPATH246.swl.thr0_state;
thread_status[985] = `IFUPATH246.swl.thr1_state;
thread_status[986] = `IFUPATH246.swl.thr2_state;
thread_status[987] = `IFUPATH246.swl.thr3_state;
thread_status[988] = `IFUPATH247.swl.thr0_state;
thread_status[989] = `IFUPATH247.swl.thr1_state;
thread_status[990] = `IFUPATH247.swl.thr2_state;
thread_status[991] = `IFUPATH247.swl.thr3_state;
thread_status[992] = `IFUPATH248.swl.thr0_state;
thread_status[993] = `IFUPATH248.swl.thr1_state;
thread_status[994] = `IFUPATH248.swl.thr2_state;
thread_status[995] = `IFUPATH248.swl.thr3_state;
thread_status[996] = `IFUPATH249.swl.thr0_state;
thread_status[997] = `IFUPATH249.swl.thr1_state;
thread_status[998] = `IFUPATH249.swl.thr2_state;
thread_status[999] = `IFUPATH249.swl.thr3_state;
thread_status[1000] = `IFUPATH250.swl.thr0_state;
thread_status[1001] = `IFUPATH250.swl.thr1_state;
thread_status[1002] = `IFUPATH250.swl.thr2_state;
thread_status[1003] = `IFUPATH250.swl.thr3_state;
thread_status[1004] = `IFUPATH251.swl.thr0_state;
thread_status[1005] = `IFUPATH251.swl.thr1_state;
thread_status[1006] = `IFUPATH251.swl.thr2_state;
thread_status[1007] = `IFUPATH251.swl.thr3_state;
thread_status[1008] = `IFUPATH252.swl.thr0_state;
thread_status[1009] = `IFUPATH252.swl.thr1_state;
thread_status[1010] = `IFUPATH252.swl.thr2_state;
thread_status[1011] = `IFUPATH252.swl.thr3_state;
thread_status[1012] = `IFUPATH253.swl.thr0_state;
thread_status[1013] = `IFUPATH253.swl.thr1_state;
thread_status[1014] = `IFUPATH253.swl.thr2_state;
thread_status[1015] = `IFUPATH253.swl.thr3_state;
thread_status[1016] = `IFUPATH254.swl.thr0_state;
thread_status[1017] = `IFUPATH254.swl.thr1_state;
thread_status[1018] = `IFUPATH254.swl.thr2_state;
thread_status[1019] = `IFUPATH254.swl.thr3_state;
thread_status[1020] = `IFUPATH255.swl.thr0_state;
thread_status[1021] = `IFUPATH255.swl.thr1_state;
thread_status[1022] = `IFUPATH255.swl.thr2_state;
thread_status[1023] = `IFUPATH255.swl.thr3_state;

    end
endtask // get_thread_status
`endif


            assign spc0_thread_id = 2'b00;
            assign spc0_rtl_pc = spc0_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(0*4)]   <= 1'b0;
                  active_thread[(0*4)+1] <= 1'b0;
                  active_thread[(0*4)+2] <= 1'b0;
                  active_thread[(0*4)+3] <= 1'b0;
                  spc0_inst_done         <= 0;
                  spc0_phy_pc_w          <= 0;
                end else begin
                  active_thread[(0*4)]   <= 1'b1;
                  active_thread[(0*4)+1] <= 1'b1;
                  active_thread[(0*4)+2] <= 1'b1;
                  active_thread[(0*4)+3] <= 1'b1;
                  spc0_inst_done         <= `TILE0.piton_pc_vld;
                  spc0_phy_pc_w          <= `TILE0.piton_pc;
                end
            end
    

            assign spc1_thread_id = 2'b00;
            assign spc1_rtl_pc = spc1_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(1*4)]   <= 1'b0;
                  active_thread[(1*4)+1] <= 1'b0;
                  active_thread[(1*4)+2] <= 1'b0;
                  active_thread[(1*4)+3] <= 1'b0;
                  spc1_inst_done         <= 0;
                  spc1_phy_pc_w          <= 0;
                end else begin
                  active_thread[(1*4)]   <= 1'b1;
                  active_thread[(1*4)+1] <= 1'b1;
                  active_thread[(1*4)+2] <= 1'b1;
                  active_thread[(1*4)+3] <= 1'b1;
                  spc1_inst_done         <= `TILE1.piton_pc_vld;
                  spc1_phy_pc_w          <= `TILE1.piton_pc;
                end
            end
    

            assign spc2_thread_id = 2'b00;
            assign spc2_rtl_pc = spc2_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(2*4)]   <= 1'b0;
                  active_thread[(2*4)+1] <= 1'b0;
                  active_thread[(2*4)+2] <= 1'b0;
                  active_thread[(2*4)+3] <= 1'b0;
                  spc2_inst_done         <= 0;
                  spc2_phy_pc_w          <= 0;
                end else begin
                  active_thread[(2*4)]   <= 1'b1;
                  active_thread[(2*4)+1] <= 1'b1;
                  active_thread[(2*4)+2] <= 1'b1;
                  active_thread[(2*4)+3] <= 1'b1;
                  spc2_inst_done         <= `TILE2.piton_pc_vld;
                  spc2_phy_pc_w          <= `TILE2.piton_pc;
                end
            end
    

            assign spc3_thread_id = 2'b00;
            assign spc3_rtl_pc = spc3_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(3*4)]   <= 1'b0;
                  active_thread[(3*4)+1] <= 1'b0;
                  active_thread[(3*4)+2] <= 1'b0;
                  active_thread[(3*4)+3] <= 1'b0;
                  spc3_inst_done         <= 0;
                  spc3_phy_pc_w          <= 0;
                end else begin
                  active_thread[(3*4)]   <= 1'b1;
                  active_thread[(3*4)+1] <= 1'b1;
                  active_thread[(3*4)+2] <= 1'b1;
                  active_thread[(3*4)+3] <= 1'b1;
                  spc3_inst_done         <= `TILE3.piton_pc_vld;
                  spc3_phy_pc_w          <= `TILE3.piton_pc;
                end
            end
    

            assign spc4_thread_id = 2'b00;
            assign spc4_rtl_pc = spc4_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(4*4)]   <= 1'b0;
                  active_thread[(4*4)+1] <= 1'b0;
                  active_thread[(4*4)+2] <= 1'b0;
                  active_thread[(4*4)+3] <= 1'b0;
                  spc4_inst_done         <= 0;
                  spc4_phy_pc_w          <= 0;
                end else begin
                  active_thread[(4*4)]   <= 1'b1;
                  active_thread[(4*4)+1] <= 1'b1;
                  active_thread[(4*4)+2] <= 1'b1;
                  active_thread[(4*4)+3] <= 1'b1;
                  spc4_inst_done         <= `TILE4.piton_pc_vld;
                  spc4_phy_pc_w          <= `TILE4.piton_pc;
                end
            end
    

            assign spc5_thread_id = 2'b00;
            assign spc5_rtl_pc = spc5_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(5*4)]   <= 1'b0;
                  active_thread[(5*4)+1] <= 1'b0;
                  active_thread[(5*4)+2] <= 1'b0;
                  active_thread[(5*4)+3] <= 1'b0;
                  spc5_inst_done         <= 0;
                  spc5_phy_pc_w          <= 0;
                end else begin
                  active_thread[(5*4)]   <= 1'b1;
                  active_thread[(5*4)+1] <= 1'b1;
                  active_thread[(5*4)+2] <= 1'b1;
                  active_thread[(5*4)+3] <= 1'b1;
                  spc5_inst_done         <= `TILE5.piton_pc_vld;
                  spc5_phy_pc_w          <= `TILE5.piton_pc;
                end
            end
    

            assign spc6_thread_id = 2'b00;
            assign spc6_rtl_pc = spc6_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(6*4)]   <= 1'b0;
                  active_thread[(6*4)+1] <= 1'b0;
                  active_thread[(6*4)+2] <= 1'b0;
                  active_thread[(6*4)+3] <= 1'b0;
                  spc6_inst_done         <= 0;
                  spc6_phy_pc_w          <= 0;
                end else begin
                  active_thread[(6*4)]   <= 1'b1;
                  active_thread[(6*4)+1] <= 1'b1;
                  active_thread[(6*4)+2] <= 1'b1;
                  active_thread[(6*4)+3] <= 1'b1;
                  spc6_inst_done         <= `TILE6.piton_pc_vld;
                  spc6_phy_pc_w          <= `TILE6.piton_pc;
                end
            end
    

            assign spc7_thread_id = 2'b00;
            assign spc7_rtl_pc = spc7_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(7*4)]   <= 1'b0;
                  active_thread[(7*4)+1] <= 1'b0;
                  active_thread[(7*4)+2] <= 1'b0;
                  active_thread[(7*4)+3] <= 1'b0;
                  spc7_inst_done         <= 0;
                  spc7_phy_pc_w          <= 0;
                end else begin
                  active_thread[(7*4)]   <= 1'b1;
                  active_thread[(7*4)+1] <= 1'b1;
                  active_thread[(7*4)+2] <= 1'b1;
                  active_thread[(7*4)+3] <= 1'b1;
                  spc7_inst_done         <= `TILE7.piton_pc_vld;
                  spc7_phy_pc_w          <= `TILE7.piton_pc;
                end
            end
    

            assign spc8_thread_id = 2'b00;
            assign spc8_rtl_pc = spc8_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(8*4)]   <= 1'b0;
                  active_thread[(8*4)+1] <= 1'b0;
                  active_thread[(8*4)+2] <= 1'b0;
                  active_thread[(8*4)+3] <= 1'b0;
                  spc8_inst_done         <= 0;
                  spc8_phy_pc_w          <= 0;
                end else begin
                  active_thread[(8*4)]   <= 1'b1;
                  active_thread[(8*4)+1] <= 1'b1;
                  active_thread[(8*4)+2] <= 1'b1;
                  active_thread[(8*4)+3] <= 1'b1;
                  spc8_inst_done         <= `TILE8.piton_pc_vld;
                  spc8_phy_pc_w          <= `TILE8.piton_pc;
                end
            end
    

            assign spc9_thread_id = 2'b00;
            assign spc9_rtl_pc = spc9_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(9*4)]   <= 1'b0;
                  active_thread[(9*4)+1] <= 1'b0;
                  active_thread[(9*4)+2] <= 1'b0;
                  active_thread[(9*4)+3] <= 1'b0;
                  spc9_inst_done         <= 0;
                  spc9_phy_pc_w          <= 0;
                end else begin
                  active_thread[(9*4)]   <= 1'b1;
                  active_thread[(9*4)+1] <= 1'b1;
                  active_thread[(9*4)+2] <= 1'b1;
                  active_thread[(9*4)+3] <= 1'b1;
                  spc9_inst_done         <= `TILE9.piton_pc_vld;
                  spc9_phy_pc_w          <= `TILE9.piton_pc;
                end
            end
    

            assign spc10_thread_id = 2'b00;
            assign spc10_rtl_pc = spc10_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(10*4)]   <= 1'b0;
                  active_thread[(10*4)+1] <= 1'b0;
                  active_thread[(10*4)+2] <= 1'b0;
                  active_thread[(10*4)+3] <= 1'b0;
                  spc10_inst_done         <= 0;
                  spc10_phy_pc_w          <= 0;
                end else begin
                  active_thread[(10*4)]   <= 1'b1;
                  active_thread[(10*4)+1] <= 1'b1;
                  active_thread[(10*4)+2] <= 1'b1;
                  active_thread[(10*4)+3] <= 1'b1;
                  spc10_inst_done         <= `TILE10.piton_pc_vld;
                  spc10_phy_pc_w          <= `TILE10.piton_pc;
                end
            end
    

            assign spc11_thread_id = 2'b00;
            assign spc11_rtl_pc = spc11_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(11*4)]   <= 1'b0;
                  active_thread[(11*4)+1] <= 1'b0;
                  active_thread[(11*4)+2] <= 1'b0;
                  active_thread[(11*4)+3] <= 1'b0;
                  spc11_inst_done         <= 0;
                  spc11_phy_pc_w          <= 0;
                end else begin
                  active_thread[(11*4)]   <= 1'b1;
                  active_thread[(11*4)+1] <= 1'b1;
                  active_thread[(11*4)+2] <= 1'b1;
                  active_thread[(11*4)+3] <= 1'b1;
                  spc11_inst_done         <= `TILE11.piton_pc_vld;
                  spc11_phy_pc_w          <= `TILE11.piton_pc;
                end
            end
    

            assign spc12_thread_id = 2'b00;
            assign spc12_rtl_pc = spc12_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(12*4)]   <= 1'b0;
                  active_thread[(12*4)+1] <= 1'b0;
                  active_thread[(12*4)+2] <= 1'b0;
                  active_thread[(12*4)+3] <= 1'b0;
                  spc12_inst_done         <= 0;
                  spc12_phy_pc_w          <= 0;
                end else begin
                  active_thread[(12*4)]   <= 1'b1;
                  active_thread[(12*4)+1] <= 1'b1;
                  active_thread[(12*4)+2] <= 1'b1;
                  active_thread[(12*4)+3] <= 1'b1;
                  spc12_inst_done         <= `TILE12.piton_pc_vld;
                  spc12_phy_pc_w          <= `TILE12.piton_pc;
                end
            end
    

            assign spc13_thread_id = 2'b00;
            assign spc13_rtl_pc = spc13_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(13*4)]   <= 1'b0;
                  active_thread[(13*4)+1] <= 1'b0;
                  active_thread[(13*4)+2] <= 1'b0;
                  active_thread[(13*4)+3] <= 1'b0;
                  spc13_inst_done         <= 0;
                  spc13_phy_pc_w          <= 0;
                end else begin
                  active_thread[(13*4)]   <= 1'b1;
                  active_thread[(13*4)+1] <= 1'b1;
                  active_thread[(13*4)+2] <= 1'b1;
                  active_thread[(13*4)+3] <= 1'b1;
                  spc13_inst_done         <= `TILE13.piton_pc_vld;
                  spc13_phy_pc_w          <= `TILE13.piton_pc;
                end
            end
    

            assign spc14_thread_id = 2'b00;
            assign spc14_rtl_pc = spc14_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(14*4)]   <= 1'b0;
                  active_thread[(14*4)+1] <= 1'b0;
                  active_thread[(14*4)+2] <= 1'b0;
                  active_thread[(14*4)+3] <= 1'b0;
                  spc14_inst_done         <= 0;
                  spc14_phy_pc_w          <= 0;
                end else begin
                  active_thread[(14*4)]   <= 1'b1;
                  active_thread[(14*4)+1] <= 1'b1;
                  active_thread[(14*4)+2] <= 1'b1;
                  active_thread[(14*4)+3] <= 1'b1;
                  spc14_inst_done         <= `TILE14.piton_pc_vld;
                  spc14_phy_pc_w          <= `TILE14.piton_pc;
                end
            end
    

            assign spc15_thread_id = 2'b00;
            assign spc15_rtl_pc = spc15_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(15*4)]   <= 1'b0;
                  active_thread[(15*4)+1] <= 1'b0;
                  active_thread[(15*4)+2] <= 1'b0;
                  active_thread[(15*4)+3] <= 1'b0;
                  spc15_inst_done         <= 0;
                  spc15_phy_pc_w          <= 0;
                end else begin
                  active_thread[(15*4)]   <= 1'b1;
                  active_thread[(15*4)+1] <= 1'b1;
                  active_thread[(15*4)+2] <= 1'b1;
                  active_thread[(15*4)+3] <= 1'b1;
                  spc15_inst_done         <= `TILE15.piton_pc_vld;
                  spc15_phy_pc_w          <= `TILE15.piton_pc;
                end
            end
    

            assign spc16_thread_id = 2'b00;
            assign spc16_rtl_pc = spc16_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(16*4)]   <= 1'b0;
                  active_thread[(16*4)+1] <= 1'b0;
                  active_thread[(16*4)+2] <= 1'b0;
                  active_thread[(16*4)+3] <= 1'b0;
                  spc16_inst_done         <= 0;
                  spc16_phy_pc_w          <= 0;
                end else begin
                  active_thread[(16*4)]   <= 1'b1;
                  active_thread[(16*4)+1] <= 1'b1;
                  active_thread[(16*4)+2] <= 1'b1;
                  active_thread[(16*4)+3] <= 1'b1;
                  spc16_inst_done         <= `TILE16.piton_pc_vld;
                  spc16_phy_pc_w          <= `TILE16.piton_pc;
                end
            end
    

            assign spc17_thread_id = 2'b00;
            assign spc17_rtl_pc = spc17_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(17*4)]   <= 1'b0;
                  active_thread[(17*4)+1] <= 1'b0;
                  active_thread[(17*4)+2] <= 1'b0;
                  active_thread[(17*4)+3] <= 1'b0;
                  spc17_inst_done         <= 0;
                  spc17_phy_pc_w          <= 0;
                end else begin
                  active_thread[(17*4)]   <= 1'b1;
                  active_thread[(17*4)+1] <= 1'b1;
                  active_thread[(17*4)+2] <= 1'b1;
                  active_thread[(17*4)+3] <= 1'b1;
                  spc17_inst_done         <= `TILE17.piton_pc_vld;
                  spc17_phy_pc_w          <= `TILE17.piton_pc;
                end
            end
    

            assign spc18_thread_id = 2'b00;
            assign spc18_rtl_pc = spc18_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(18*4)]   <= 1'b0;
                  active_thread[(18*4)+1] <= 1'b0;
                  active_thread[(18*4)+2] <= 1'b0;
                  active_thread[(18*4)+3] <= 1'b0;
                  spc18_inst_done         <= 0;
                  spc18_phy_pc_w          <= 0;
                end else begin
                  active_thread[(18*4)]   <= 1'b1;
                  active_thread[(18*4)+1] <= 1'b1;
                  active_thread[(18*4)+2] <= 1'b1;
                  active_thread[(18*4)+3] <= 1'b1;
                  spc18_inst_done         <= `TILE18.piton_pc_vld;
                  spc18_phy_pc_w          <= `TILE18.piton_pc;
                end
            end
    

            assign spc19_thread_id = 2'b00;
            assign spc19_rtl_pc = spc19_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(19*4)]   <= 1'b0;
                  active_thread[(19*4)+1] <= 1'b0;
                  active_thread[(19*4)+2] <= 1'b0;
                  active_thread[(19*4)+3] <= 1'b0;
                  spc19_inst_done         <= 0;
                  spc19_phy_pc_w          <= 0;
                end else begin
                  active_thread[(19*4)]   <= 1'b1;
                  active_thread[(19*4)+1] <= 1'b1;
                  active_thread[(19*4)+2] <= 1'b1;
                  active_thread[(19*4)+3] <= 1'b1;
                  spc19_inst_done         <= `TILE19.piton_pc_vld;
                  spc19_phy_pc_w          <= `TILE19.piton_pc;
                end
            end
    

            assign spc20_thread_id = 2'b00;
            assign spc20_rtl_pc = spc20_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(20*4)]   <= 1'b0;
                  active_thread[(20*4)+1] <= 1'b0;
                  active_thread[(20*4)+2] <= 1'b0;
                  active_thread[(20*4)+3] <= 1'b0;
                  spc20_inst_done         <= 0;
                  spc20_phy_pc_w          <= 0;
                end else begin
                  active_thread[(20*4)]   <= 1'b1;
                  active_thread[(20*4)+1] <= 1'b1;
                  active_thread[(20*4)+2] <= 1'b1;
                  active_thread[(20*4)+3] <= 1'b1;
                  spc20_inst_done         <= `TILE20.piton_pc_vld;
                  spc20_phy_pc_w          <= `TILE20.piton_pc;
                end
            end
    

            assign spc21_thread_id = 2'b00;
            assign spc21_rtl_pc = spc21_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(21*4)]   <= 1'b0;
                  active_thread[(21*4)+1] <= 1'b0;
                  active_thread[(21*4)+2] <= 1'b0;
                  active_thread[(21*4)+3] <= 1'b0;
                  spc21_inst_done         <= 0;
                  spc21_phy_pc_w          <= 0;
                end else begin
                  active_thread[(21*4)]   <= 1'b1;
                  active_thread[(21*4)+1] <= 1'b1;
                  active_thread[(21*4)+2] <= 1'b1;
                  active_thread[(21*4)+3] <= 1'b1;
                  spc21_inst_done         <= `TILE21.piton_pc_vld;
                  spc21_phy_pc_w          <= `TILE21.piton_pc;
                end
            end
    

            assign spc22_thread_id = 2'b00;
            assign spc22_rtl_pc = spc22_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(22*4)]   <= 1'b0;
                  active_thread[(22*4)+1] <= 1'b0;
                  active_thread[(22*4)+2] <= 1'b0;
                  active_thread[(22*4)+3] <= 1'b0;
                  spc22_inst_done         <= 0;
                  spc22_phy_pc_w          <= 0;
                end else begin
                  active_thread[(22*4)]   <= 1'b1;
                  active_thread[(22*4)+1] <= 1'b1;
                  active_thread[(22*4)+2] <= 1'b1;
                  active_thread[(22*4)+3] <= 1'b1;
                  spc22_inst_done         <= `TILE22.piton_pc_vld;
                  spc22_phy_pc_w          <= `TILE22.piton_pc;
                end
            end
    

            assign spc23_thread_id = 2'b00;
            assign spc23_rtl_pc = spc23_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(23*4)]   <= 1'b0;
                  active_thread[(23*4)+1] <= 1'b0;
                  active_thread[(23*4)+2] <= 1'b0;
                  active_thread[(23*4)+3] <= 1'b0;
                  spc23_inst_done         <= 0;
                  spc23_phy_pc_w          <= 0;
                end else begin
                  active_thread[(23*4)]   <= 1'b1;
                  active_thread[(23*4)+1] <= 1'b1;
                  active_thread[(23*4)+2] <= 1'b1;
                  active_thread[(23*4)+3] <= 1'b1;
                  spc23_inst_done         <= `TILE23.piton_pc_vld;
                  spc23_phy_pc_w          <= `TILE23.piton_pc;
                end
            end
    

            assign spc24_thread_id = 2'b00;
            assign spc24_rtl_pc = spc24_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(24*4)]   <= 1'b0;
                  active_thread[(24*4)+1] <= 1'b0;
                  active_thread[(24*4)+2] <= 1'b0;
                  active_thread[(24*4)+3] <= 1'b0;
                  spc24_inst_done         <= 0;
                  spc24_phy_pc_w          <= 0;
                end else begin
                  active_thread[(24*4)]   <= 1'b1;
                  active_thread[(24*4)+1] <= 1'b1;
                  active_thread[(24*4)+2] <= 1'b1;
                  active_thread[(24*4)+3] <= 1'b1;
                  spc24_inst_done         <= `TILE24.piton_pc_vld;
                  spc24_phy_pc_w          <= `TILE24.piton_pc;
                end
            end
    

            assign spc25_thread_id = 2'b00;
            assign spc25_rtl_pc = spc25_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(25*4)]   <= 1'b0;
                  active_thread[(25*4)+1] <= 1'b0;
                  active_thread[(25*4)+2] <= 1'b0;
                  active_thread[(25*4)+3] <= 1'b0;
                  spc25_inst_done         <= 0;
                  spc25_phy_pc_w          <= 0;
                end else begin
                  active_thread[(25*4)]   <= 1'b1;
                  active_thread[(25*4)+1] <= 1'b1;
                  active_thread[(25*4)+2] <= 1'b1;
                  active_thread[(25*4)+3] <= 1'b1;
                  spc25_inst_done         <= `TILE25.piton_pc_vld;
                  spc25_phy_pc_w          <= `TILE25.piton_pc;
                end
            end
    

            assign spc26_thread_id = 2'b00;
            assign spc26_rtl_pc = spc26_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(26*4)]   <= 1'b0;
                  active_thread[(26*4)+1] <= 1'b0;
                  active_thread[(26*4)+2] <= 1'b0;
                  active_thread[(26*4)+3] <= 1'b0;
                  spc26_inst_done         <= 0;
                  spc26_phy_pc_w          <= 0;
                end else begin
                  active_thread[(26*4)]   <= 1'b1;
                  active_thread[(26*4)+1] <= 1'b1;
                  active_thread[(26*4)+2] <= 1'b1;
                  active_thread[(26*4)+3] <= 1'b1;
                  spc26_inst_done         <= `TILE26.piton_pc_vld;
                  spc26_phy_pc_w          <= `TILE26.piton_pc;
                end
            end
    

            assign spc27_thread_id = 2'b00;
            assign spc27_rtl_pc = spc27_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(27*4)]   <= 1'b0;
                  active_thread[(27*4)+1] <= 1'b0;
                  active_thread[(27*4)+2] <= 1'b0;
                  active_thread[(27*4)+3] <= 1'b0;
                  spc27_inst_done         <= 0;
                  spc27_phy_pc_w          <= 0;
                end else begin
                  active_thread[(27*4)]   <= 1'b1;
                  active_thread[(27*4)+1] <= 1'b1;
                  active_thread[(27*4)+2] <= 1'b1;
                  active_thread[(27*4)+3] <= 1'b1;
                  spc27_inst_done         <= `TILE27.piton_pc_vld;
                  spc27_phy_pc_w          <= `TILE27.piton_pc;
                end
            end
    

            assign spc28_thread_id = 2'b00;
            assign spc28_rtl_pc = spc28_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(28*4)]   <= 1'b0;
                  active_thread[(28*4)+1] <= 1'b0;
                  active_thread[(28*4)+2] <= 1'b0;
                  active_thread[(28*4)+3] <= 1'b0;
                  spc28_inst_done         <= 0;
                  spc28_phy_pc_w          <= 0;
                end else begin
                  active_thread[(28*4)]   <= 1'b1;
                  active_thread[(28*4)+1] <= 1'b1;
                  active_thread[(28*4)+2] <= 1'b1;
                  active_thread[(28*4)+3] <= 1'b1;
                  spc28_inst_done         <= `TILE28.piton_pc_vld;
                  spc28_phy_pc_w          <= `TILE28.piton_pc;
                end
            end
    

            assign spc29_thread_id = 2'b00;
            assign spc29_rtl_pc = spc29_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(29*4)]   <= 1'b0;
                  active_thread[(29*4)+1] <= 1'b0;
                  active_thread[(29*4)+2] <= 1'b0;
                  active_thread[(29*4)+3] <= 1'b0;
                  spc29_inst_done         <= 0;
                  spc29_phy_pc_w          <= 0;
                end else begin
                  active_thread[(29*4)]   <= 1'b1;
                  active_thread[(29*4)+1] <= 1'b1;
                  active_thread[(29*4)+2] <= 1'b1;
                  active_thread[(29*4)+3] <= 1'b1;
                  spc29_inst_done         <= `TILE29.piton_pc_vld;
                  spc29_phy_pc_w          <= `TILE29.piton_pc;
                end
            end
    

            assign spc30_thread_id = 2'b00;
            assign spc30_rtl_pc = spc30_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(30*4)]   <= 1'b0;
                  active_thread[(30*4)+1] <= 1'b0;
                  active_thread[(30*4)+2] <= 1'b0;
                  active_thread[(30*4)+3] <= 1'b0;
                  spc30_inst_done         <= 0;
                  spc30_phy_pc_w          <= 0;
                end else begin
                  active_thread[(30*4)]   <= 1'b1;
                  active_thread[(30*4)+1] <= 1'b1;
                  active_thread[(30*4)+2] <= 1'b1;
                  active_thread[(30*4)+3] <= 1'b1;
                  spc30_inst_done         <= `TILE30.piton_pc_vld;
                  spc30_phy_pc_w          <= `TILE30.piton_pc;
                end
            end
    

            assign spc31_thread_id = 2'b00;
            assign spc31_rtl_pc = spc31_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(31*4)]   <= 1'b0;
                  active_thread[(31*4)+1] <= 1'b0;
                  active_thread[(31*4)+2] <= 1'b0;
                  active_thread[(31*4)+3] <= 1'b0;
                  spc31_inst_done         <= 0;
                  spc31_phy_pc_w          <= 0;
                end else begin
                  active_thread[(31*4)]   <= 1'b1;
                  active_thread[(31*4)+1] <= 1'b1;
                  active_thread[(31*4)+2] <= 1'b1;
                  active_thread[(31*4)+3] <= 1'b1;
                  spc31_inst_done         <= `TILE31.piton_pc_vld;
                  spc31_phy_pc_w          <= `TILE31.piton_pc;
                end
            end
    

            assign spc32_thread_id = 2'b00;
            assign spc32_rtl_pc = spc32_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(32*4)]   <= 1'b0;
                  active_thread[(32*4)+1] <= 1'b0;
                  active_thread[(32*4)+2] <= 1'b0;
                  active_thread[(32*4)+3] <= 1'b0;
                  spc32_inst_done         <= 0;
                  spc32_phy_pc_w          <= 0;
                end else begin
                  active_thread[(32*4)]   <= 1'b1;
                  active_thread[(32*4)+1] <= 1'b1;
                  active_thread[(32*4)+2] <= 1'b1;
                  active_thread[(32*4)+3] <= 1'b1;
                  spc32_inst_done         <= `TILE32.piton_pc_vld;
                  spc32_phy_pc_w          <= `TILE32.piton_pc;
                end
            end
    

            assign spc33_thread_id = 2'b00;
            assign spc33_rtl_pc = spc33_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(33*4)]   <= 1'b0;
                  active_thread[(33*4)+1] <= 1'b0;
                  active_thread[(33*4)+2] <= 1'b0;
                  active_thread[(33*4)+3] <= 1'b0;
                  spc33_inst_done         <= 0;
                  spc33_phy_pc_w          <= 0;
                end else begin
                  active_thread[(33*4)]   <= 1'b1;
                  active_thread[(33*4)+1] <= 1'b1;
                  active_thread[(33*4)+2] <= 1'b1;
                  active_thread[(33*4)+3] <= 1'b1;
                  spc33_inst_done         <= `TILE33.piton_pc_vld;
                  spc33_phy_pc_w          <= `TILE33.piton_pc;
                end
            end
    

            assign spc34_thread_id = 2'b00;
            assign spc34_rtl_pc = spc34_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(34*4)]   <= 1'b0;
                  active_thread[(34*4)+1] <= 1'b0;
                  active_thread[(34*4)+2] <= 1'b0;
                  active_thread[(34*4)+3] <= 1'b0;
                  spc34_inst_done         <= 0;
                  spc34_phy_pc_w          <= 0;
                end else begin
                  active_thread[(34*4)]   <= 1'b1;
                  active_thread[(34*4)+1] <= 1'b1;
                  active_thread[(34*4)+2] <= 1'b1;
                  active_thread[(34*4)+3] <= 1'b1;
                  spc34_inst_done         <= `TILE34.piton_pc_vld;
                  spc34_phy_pc_w          <= `TILE34.piton_pc;
                end
            end
    

            assign spc35_thread_id = 2'b00;
            assign spc35_rtl_pc = spc35_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(35*4)]   <= 1'b0;
                  active_thread[(35*4)+1] <= 1'b0;
                  active_thread[(35*4)+2] <= 1'b0;
                  active_thread[(35*4)+3] <= 1'b0;
                  spc35_inst_done         <= 0;
                  spc35_phy_pc_w          <= 0;
                end else begin
                  active_thread[(35*4)]   <= 1'b1;
                  active_thread[(35*4)+1] <= 1'b1;
                  active_thread[(35*4)+2] <= 1'b1;
                  active_thread[(35*4)+3] <= 1'b1;
                  spc35_inst_done         <= `TILE35.piton_pc_vld;
                  spc35_phy_pc_w          <= `TILE35.piton_pc;
                end
            end
    

            assign spc36_thread_id = 2'b00;
            assign spc36_rtl_pc = spc36_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(36*4)]   <= 1'b0;
                  active_thread[(36*4)+1] <= 1'b0;
                  active_thread[(36*4)+2] <= 1'b0;
                  active_thread[(36*4)+3] <= 1'b0;
                  spc36_inst_done         <= 0;
                  spc36_phy_pc_w          <= 0;
                end else begin
                  active_thread[(36*4)]   <= 1'b1;
                  active_thread[(36*4)+1] <= 1'b1;
                  active_thread[(36*4)+2] <= 1'b1;
                  active_thread[(36*4)+3] <= 1'b1;
                  spc36_inst_done         <= `TILE36.piton_pc_vld;
                  spc36_phy_pc_w          <= `TILE36.piton_pc;
                end
            end
    

            assign spc37_thread_id = 2'b00;
            assign spc37_rtl_pc = spc37_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(37*4)]   <= 1'b0;
                  active_thread[(37*4)+1] <= 1'b0;
                  active_thread[(37*4)+2] <= 1'b0;
                  active_thread[(37*4)+3] <= 1'b0;
                  spc37_inst_done         <= 0;
                  spc37_phy_pc_w          <= 0;
                end else begin
                  active_thread[(37*4)]   <= 1'b1;
                  active_thread[(37*4)+1] <= 1'b1;
                  active_thread[(37*4)+2] <= 1'b1;
                  active_thread[(37*4)+3] <= 1'b1;
                  spc37_inst_done         <= `TILE37.piton_pc_vld;
                  spc37_phy_pc_w          <= `TILE37.piton_pc;
                end
            end
    

            assign spc38_thread_id = 2'b00;
            assign spc38_rtl_pc = spc38_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(38*4)]   <= 1'b0;
                  active_thread[(38*4)+1] <= 1'b0;
                  active_thread[(38*4)+2] <= 1'b0;
                  active_thread[(38*4)+3] <= 1'b0;
                  spc38_inst_done         <= 0;
                  spc38_phy_pc_w          <= 0;
                end else begin
                  active_thread[(38*4)]   <= 1'b1;
                  active_thread[(38*4)+1] <= 1'b1;
                  active_thread[(38*4)+2] <= 1'b1;
                  active_thread[(38*4)+3] <= 1'b1;
                  spc38_inst_done         <= `TILE38.piton_pc_vld;
                  spc38_phy_pc_w          <= `TILE38.piton_pc;
                end
            end
    

            assign spc39_thread_id = 2'b00;
            assign spc39_rtl_pc = spc39_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(39*4)]   <= 1'b0;
                  active_thread[(39*4)+1] <= 1'b0;
                  active_thread[(39*4)+2] <= 1'b0;
                  active_thread[(39*4)+3] <= 1'b0;
                  spc39_inst_done         <= 0;
                  spc39_phy_pc_w          <= 0;
                end else begin
                  active_thread[(39*4)]   <= 1'b1;
                  active_thread[(39*4)+1] <= 1'b1;
                  active_thread[(39*4)+2] <= 1'b1;
                  active_thread[(39*4)+3] <= 1'b1;
                  spc39_inst_done         <= `TILE39.piton_pc_vld;
                  spc39_phy_pc_w          <= `TILE39.piton_pc;
                end
            end
    

            assign spc40_thread_id = 2'b00;
            assign spc40_rtl_pc = spc40_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(40*4)]   <= 1'b0;
                  active_thread[(40*4)+1] <= 1'b0;
                  active_thread[(40*4)+2] <= 1'b0;
                  active_thread[(40*4)+3] <= 1'b0;
                  spc40_inst_done         <= 0;
                  spc40_phy_pc_w          <= 0;
                end else begin
                  active_thread[(40*4)]   <= 1'b1;
                  active_thread[(40*4)+1] <= 1'b1;
                  active_thread[(40*4)+2] <= 1'b1;
                  active_thread[(40*4)+3] <= 1'b1;
                  spc40_inst_done         <= `TILE40.piton_pc_vld;
                  spc40_phy_pc_w          <= `TILE40.piton_pc;
                end
            end
    

            assign spc41_thread_id = 2'b00;
            assign spc41_rtl_pc = spc41_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(41*4)]   <= 1'b0;
                  active_thread[(41*4)+1] <= 1'b0;
                  active_thread[(41*4)+2] <= 1'b0;
                  active_thread[(41*4)+3] <= 1'b0;
                  spc41_inst_done         <= 0;
                  spc41_phy_pc_w          <= 0;
                end else begin
                  active_thread[(41*4)]   <= 1'b1;
                  active_thread[(41*4)+1] <= 1'b1;
                  active_thread[(41*4)+2] <= 1'b1;
                  active_thread[(41*4)+3] <= 1'b1;
                  spc41_inst_done         <= `TILE41.piton_pc_vld;
                  spc41_phy_pc_w          <= `TILE41.piton_pc;
                end
            end
    

            assign spc42_thread_id = 2'b00;
            assign spc42_rtl_pc = spc42_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(42*4)]   <= 1'b0;
                  active_thread[(42*4)+1] <= 1'b0;
                  active_thread[(42*4)+2] <= 1'b0;
                  active_thread[(42*4)+3] <= 1'b0;
                  spc42_inst_done         <= 0;
                  spc42_phy_pc_w          <= 0;
                end else begin
                  active_thread[(42*4)]   <= 1'b1;
                  active_thread[(42*4)+1] <= 1'b1;
                  active_thread[(42*4)+2] <= 1'b1;
                  active_thread[(42*4)+3] <= 1'b1;
                  spc42_inst_done         <= `TILE42.piton_pc_vld;
                  spc42_phy_pc_w          <= `TILE42.piton_pc;
                end
            end
    

            assign spc43_thread_id = 2'b00;
            assign spc43_rtl_pc = spc43_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(43*4)]   <= 1'b0;
                  active_thread[(43*4)+1] <= 1'b0;
                  active_thread[(43*4)+2] <= 1'b0;
                  active_thread[(43*4)+3] <= 1'b0;
                  spc43_inst_done         <= 0;
                  spc43_phy_pc_w          <= 0;
                end else begin
                  active_thread[(43*4)]   <= 1'b1;
                  active_thread[(43*4)+1] <= 1'b1;
                  active_thread[(43*4)+2] <= 1'b1;
                  active_thread[(43*4)+3] <= 1'b1;
                  spc43_inst_done         <= `TILE43.piton_pc_vld;
                  spc43_phy_pc_w          <= `TILE43.piton_pc;
                end
            end
    

            assign spc44_thread_id = 2'b00;
            assign spc44_rtl_pc = spc44_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(44*4)]   <= 1'b0;
                  active_thread[(44*4)+1] <= 1'b0;
                  active_thread[(44*4)+2] <= 1'b0;
                  active_thread[(44*4)+3] <= 1'b0;
                  spc44_inst_done         <= 0;
                  spc44_phy_pc_w          <= 0;
                end else begin
                  active_thread[(44*4)]   <= 1'b1;
                  active_thread[(44*4)+1] <= 1'b1;
                  active_thread[(44*4)+2] <= 1'b1;
                  active_thread[(44*4)+3] <= 1'b1;
                  spc44_inst_done         <= `TILE44.piton_pc_vld;
                  spc44_phy_pc_w          <= `TILE44.piton_pc;
                end
            end
    

            assign spc45_thread_id = 2'b00;
            assign spc45_rtl_pc = spc45_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(45*4)]   <= 1'b0;
                  active_thread[(45*4)+1] <= 1'b0;
                  active_thread[(45*4)+2] <= 1'b0;
                  active_thread[(45*4)+3] <= 1'b0;
                  spc45_inst_done         <= 0;
                  spc45_phy_pc_w          <= 0;
                end else begin
                  active_thread[(45*4)]   <= 1'b1;
                  active_thread[(45*4)+1] <= 1'b1;
                  active_thread[(45*4)+2] <= 1'b1;
                  active_thread[(45*4)+3] <= 1'b1;
                  spc45_inst_done         <= `TILE45.piton_pc_vld;
                  spc45_phy_pc_w          <= `TILE45.piton_pc;
                end
            end
    

            assign spc46_thread_id = 2'b00;
            assign spc46_rtl_pc = spc46_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(46*4)]   <= 1'b0;
                  active_thread[(46*4)+1] <= 1'b0;
                  active_thread[(46*4)+2] <= 1'b0;
                  active_thread[(46*4)+3] <= 1'b0;
                  spc46_inst_done         <= 0;
                  spc46_phy_pc_w          <= 0;
                end else begin
                  active_thread[(46*4)]   <= 1'b1;
                  active_thread[(46*4)+1] <= 1'b1;
                  active_thread[(46*4)+2] <= 1'b1;
                  active_thread[(46*4)+3] <= 1'b1;
                  spc46_inst_done         <= `TILE46.piton_pc_vld;
                  spc46_phy_pc_w          <= `TILE46.piton_pc;
                end
            end
    

            assign spc47_thread_id = 2'b00;
            assign spc47_rtl_pc = spc47_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(47*4)]   <= 1'b0;
                  active_thread[(47*4)+1] <= 1'b0;
                  active_thread[(47*4)+2] <= 1'b0;
                  active_thread[(47*4)+3] <= 1'b0;
                  spc47_inst_done         <= 0;
                  spc47_phy_pc_w          <= 0;
                end else begin
                  active_thread[(47*4)]   <= 1'b1;
                  active_thread[(47*4)+1] <= 1'b1;
                  active_thread[(47*4)+2] <= 1'b1;
                  active_thread[(47*4)+3] <= 1'b1;
                  spc47_inst_done         <= `TILE47.piton_pc_vld;
                  spc47_phy_pc_w          <= `TILE47.piton_pc;
                end
            end
    

            assign spc48_thread_id = 2'b00;
            assign spc48_rtl_pc = spc48_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(48*4)]   <= 1'b0;
                  active_thread[(48*4)+1] <= 1'b0;
                  active_thread[(48*4)+2] <= 1'b0;
                  active_thread[(48*4)+3] <= 1'b0;
                  spc48_inst_done         <= 0;
                  spc48_phy_pc_w          <= 0;
                end else begin
                  active_thread[(48*4)]   <= 1'b1;
                  active_thread[(48*4)+1] <= 1'b1;
                  active_thread[(48*4)+2] <= 1'b1;
                  active_thread[(48*4)+3] <= 1'b1;
                  spc48_inst_done         <= `TILE48.piton_pc_vld;
                  spc48_phy_pc_w          <= `TILE48.piton_pc;
                end
            end
    

            assign spc49_thread_id = 2'b00;
            assign spc49_rtl_pc = spc49_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(49*4)]   <= 1'b0;
                  active_thread[(49*4)+1] <= 1'b0;
                  active_thread[(49*4)+2] <= 1'b0;
                  active_thread[(49*4)+3] <= 1'b0;
                  spc49_inst_done         <= 0;
                  spc49_phy_pc_w          <= 0;
                end else begin
                  active_thread[(49*4)]   <= 1'b1;
                  active_thread[(49*4)+1] <= 1'b1;
                  active_thread[(49*4)+2] <= 1'b1;
                  active_thread[(49*4)+3] <= 1'b1;
                  spc49_inst_done         <= `TILE49.piton_pc_vld;
                  spc49_phy_pc_w          <= `TILE49.piton_pc;
                end
            end
    

            assign spc50_thread_id = 2'b00;
            assign spc50_rtl_pc = spc50_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(50*4)]   <= 1'b0;
                  active_thread[(50*4)+1] <= 1'b0;
                  active_thread[(50*4)+2] <= 1'b0;
                  active_thread[(50*4)+3] <= 1'b0;
                  spc50_inst_done         <= 0;
                  spc50_phy_pc_w          <= 0;
                end else begin
                  active_thread[(50*4)]   <= 1'b1;
                  active_thread[(50*4)+1] <= 1'b1;
                  active_thread[(50*4)+2] <= 1'b1;
                  active_thread[(50*4)+3] <= 1'b1;
                  spc50_inst_done         <= `TILE50.piton_pc_vld;
                  spc50_phy_pc_w          <= `TILE50.piton_pc;
                end
            end
    

            assign spc51_thread_id = 2'b00;
            assign spc51_rtl_pc = spc51_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(51*4)]   <= 1'b0;
                  active_thread[(51*4)+1] <= 1'b0;
                  active_thread[(51*4)+2] <= 1'b0;
                  active_thread[(51*4)+3] <= 1'b0;
                  spc51_inst_done         <= 0;
                  spc51_phy_pc_w          <= 0;
                end else begin
                  active_thread[(51*4)]   <= 1'b1;
                  active_thread[(51*4)+1] <= 1'b1;
                  active_thread[(51*4)+2] <= 1'b1;
                  active_thread[(51*4)+3] <= 1'b1;
                  spc51_inst_done         <= `TILE51.piton_pc_vld;
                  spc51_phy_pc_w          <= `TILE51.piton_pc;
                end
            end
    

            assign spc52_thread_id = 2'b00;
            assign spc52_rtl_pc = spc52_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(52*4)]   <= 1'b0;
                  active_thread[(52*4)+1] <= 1'b0;
                  active_thread[(52*4)+2] <= 1'b0;
                  active_thread[(52*4)+3] <= 1'b0;
                  spc52_inst_done         <= 0;
                  spc52_phy_pc_w          <= 0;
                end else begin
                  active_thread[(52*4)]   <= 1'b1;
                  active_thread[(52*4)+1] <= 1'b1;
                  active_thread[(52*4)+2] <= 1'b1;
                  active_thread[(52*4)+3] <= 1'b1;
                  spc52_inst_done         <= `TILE52.piton_pc_vld;
                  spc52_phy_pc_w          <= `TILE52.piton_pc;
                end
            end
    

            assign spc53_thread_id = 2'b00;
            assign spc53_rtl_pc = spc53_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(53*4)]   <= 1'b0;
                  active_thread[(53*4)+1] <= 1'b0;
                  active_thread[(53*4)+2] <= 1'b0;
                  active_thread[(53*4)+3] <= 1'b0;
                  spc53_inst_done         <= 0;
                  spc53_phy_pc_w          <= 0;
                end else begin
                  active_thread[(53*4)]   <= 1'b1;
                  active_thread[(53*4)+1] <= 1'b1;
                  active_thread[(53*4)+2] <= 1'b1;
                  active_thread[(53*4)+3] <= 1'b1;
                  spc53_inst_done         <= `TILE53.piton_pc_vld;
                  spc53_phy_pc_w          <= `TILE53.piton_pc;
                end
            end
    

            assign spc54_thread_id = 2'b00;
            assign spc54_rtl_pc = spc54_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(54*4)]   <= 1'b0;
                  active_thread[(54*4)+1] <= 1'b0;
                  active_thread[(54*4)+2] <= 1'b0;
                  active_thread[(54*4)+3] <= 1'b0;
                  spc54_inst_done         <= 0;
                  spc54_phy_pc_w          <= 0;
                end else begin
                  active_thread[(54*4)]   <= 1'b1;
                  active_thread[(54*4)+1] <= 1'b1;
                  active_thread[(54*4)+2] <= 1'b1;
                  active_thread[(54*4)+3] <= 1'b1;
                  spc54_inst_done         <= `TILE54.piton_pc_vld;
                  spc54_phy_pc_w          <= `TILE54.piton_pc;
                end
            end
    

            assign spc55_thread_id = 2'b00;
            assign spc55_rtl_pc = spc55_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(55*4)]   <= 1'b0;
                  active_thread[(55*4)+1] <= 1'b0;
                  active_thread[(55*4)+2] <= 1'b0;
                  active_thread[(55*4)+3] <= 1'b0;
                  spc55_inst_done         <= 0;
                  spc55_phy_pc_w          <= 0;
                end else begin
                  active_thread[(55*4)]   <= 1'b1;
                  active_thread[(55*4)+1] <= 1'b1;
                  active_thread[(55*4)+2] <= 1'b1;
                  active_thread[(55*4)+3] <= 1'b1;
                  spc55_inst_done         <= `TILE55.piton_pc_vld;
                  spc55_phy_pc_w          <= `TILE55.piton_pc;
                end
            end
    

            assign spc56_thread_id = 2'b00;
            assign spc56_rtl_pc = spc56_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(56*4)]   <= 1'b0;
                  active_thread[(56*4)+1] <= 1'b0;
                  active_thread[(56*4)+2] <= 1'b0;
                  active_thread[(56*4)+3] <= 1'b0;
                  spc56_inst_done         <= 0;
                  spc56_phy_pc_w          <= 0;
                end else begin
                  active_thread[(56*4)]   <= 1'b1;
                  active_thread[(56*4)+1] <= 1'b1;
                  active_thread[(56*4)+2] <= 1'b1;
                  active_thread[(56*4)+3] <= 1'b1;
                  spc56_inst_done         <= `TILE56.piton_pc_vld;
                  spc56_phy_pc_w          <= `TILE56.piton_pc;
                end
            end
    

            assign spc57_thread_id = 2'b00;
            assign spc57_rtl_pc = spc57_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(57*4)]   <= 1'b0;
                  active_thread[(57*4)+1] <= 1'b0;
                  active_thread[(57*4)+2] <= 1'b0;
                  active_thread[(57*4)+3] <= 1'b0;
                  spc57_inst_done         <= 0;
                  spc57_phy_pc_w          <= 0;
                end else begin
                  active_thread[(57*4)]   <= 1'b1;
                  active_thread[(57*4)+1] <= 1'b1;
                  active_thread[(57*4)+2] <= 1'b1;
                  active_thread[(57*4)+3] <= 1'b1;
                  spc57_inst_done         <= `TILE57.piton_pc_vld;
                  spc57_phy_pc_w          <= `TILE57.piton_pc;
                end
            end
    

            assign spc58_thread_id = 2'b00;
            assign spc58_rtl_pc = spc58_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(58*4)]   <= 1'b0;
                  active_thread[(58*4)+1] <= 1'b0;
                  active_thread[(58*4)+2] <= 1'b0;
                  active_thread[(58*4)+3] <= 1'b0;
                  spc58_inst_done         <= 0;
                  spc58_phy_pc_w          <= 0;
                end else begin
                  active_thread[(58*4)]   <= 1'b1;
                  active_thread[(58*4)+1] <= 1'b1;
                  active_thread[(58*4)+2] <= 1'b1;
                  active_thread[(58*4)+3] <= 1'b1;
                  spc58_inst_done         <= `TILE58.piton_pc_vld;
                  spc58_phy_pc_w          <= `TILE58.piton_pc;
                end
            end
    

            assign spc59_thread_id = 2'b00;
            assign spc59_rtl_pc = spc59_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(59*4)]   <= 1'b0;
                  active_thread[(59*4)+1] <= 1'b0;
                  active_thread[(59*4)+2] <= 1'b0;
                  active_thread[(59*4)+3] <= 1'b0;
                  spc59_inst_done         <= 0;
                  spc59_phy_pc_w          <= 0;
                end else begin
                  active_thread[(59*4)]   <= 1'b1;
                  active_thread[(59*4)+1] <= 1'b1;
                  active_thread[(59*4)+2] <= 1'b1;
                  active_thread[(59*4)+3] <= 1'b1;
                  spc59_inst_done         <= `TILE59.piton_pc_vld;
                  spc59_phy_pc_w          <= `TILE59.piton_pc;
                end
            end
    

            assign spc60_thread_id = 2'b00;
            assign spc60_rtl_pc = spc60_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(60*4)]   <= 1'b0;
                  active_thread[(60*4)+1] <= 1'b0;
                  active_thread[(60*4)+2] <= 1'b0;
                  active_thread[(60*4)+3] <= 1'b0;
                  spc60_inst_done         <= 0;
                  spc60_phy_pc_w          <= 0;
                end else begin
                  active_thread[(60*4)]   <= 1'b1;
                  active_thread[(60*4)+1] <= 1'b1;
                  active_thread[(60*4)+2] <= 1'b1;
                  active_thread[(60*4)+3] <= 1'b1;
                  spc60_inst_done         <= `TILE60.piton_pc_vld;
                  spc60_phy_pc_w          <= `TILE60.piton_pc;
                end
            end
    

            assign spc61_thread_id = 2'b00;
            assign spc61_rtl_pc = spc61_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(61*4)]   <= 1'b0;
                  active_thread[(61*4)+1] <= 1'b0;
                  active_thread[(61*4)+2] <= 1'b0;
                  active_thread[(61*4)+3] <= 1'b0;
                  spc61_inst_done         <= 0;
                  spc61_phy_pc_w          <= 0;
                end else begin
                  active_thread[(61*4)]   <= 1'b1;
                  active_thread[(61*4)+1] <= 1'b1;
                  active_thread[(61*4)+2] <= 1'b1;
                  active_thread[(61*4)+3] <= 1'b1;
                  spc61_inst_done         <= `TILE61.piton_pc_vld;
                  spc61_phy_pc_w          <= `TILE61.piton_pc;
                end
            end
    

            assign spc62_thread_id = 2'b00;
            assign spc62_rtl_pc = spc62_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(62*4)]   <= 1'b0;
                  active_thread[(62*4)+1] <= 1'b0;
                  active_thread[(62*4)+2] <= 1'b0;
                  active_thread[(62*4)+3] <= 1'b0;
                  spc62_inst_done         <= 0;
                  spc62_phy_pc_w          <= 0;
                end else begin
                  active_thread[(62*4)]   <= 1'b1;
                  active_thread[(62*4)+1] <= 1'b1;
                  active_thread[(62*4)+2] <= 1'b1;
                  active_thread[(62*4)+3] <= 1'b1;
                  spc62_inst_done         <= `TILE62.piton_pc_vld;
                  spc62_phy_pc_w          <= `TILE62.piton_pc;
                end
            end
    

            assign spc63_thread_id = 2'b00;
            assign spc63_rtl_pc = spc63_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(63*4)]   <= 1'b0;
                  active_thread[(63*4)+1] <= 1'b0;
                  active_thread[(63*4)+2] <= 1'b0;
                  active_thread[(63*4)+3] <= 1'b0;
                  spc63_inst_done         <= 0;
                  spc63_phy_pc_w          <= 0;
                end else begin
                  active_thread[(63*4)]   <= 1'b1;
                  active_thread[(63*4)+1] <= 1'b1;
                  active_thread[(63*4)+2] <= 1'b1;
                  active_thread[(63*4)+3] <= 1'b1;
                  spc63_inst_done         <= `TILE63.piton_pc_vld;
                  spc63_phy_pc_w          <= `TILE63.piton_pc;
                end
            end
    

            assign spc64_thread_id = 2'b00;
            assign spc64_rtl_pc = spc64_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(64*4)]   <= 1'b0;
                  active_thread[(64*4)+1] <= 1'b0;
                  active_thread[(64*4)+2] <= 1'b0;
                  active_thread[(64*4)+3] <= 1'b0;
                  spc64_inst_done         <= 0;
                  spc64_phy_pc_w          <= 0;
                end else begin
                  active_thread[(64*4)]   <= 1'b1;
                  active_thread[(64*4)+1] <= 1'b1;
                  active_thread[(64*4)+2] <= 1'b1;
                  active_thread[(64*4)+3] <= 1'b1;
                  spc64_inst_done         <= `TILE64.piton_pc_vld;
                  spc64_phy_pc_w          <= `TILE64.piton_pc;
                end
            end
    

            assign spc65_thread_id = 2'b00;
            assign spc65_rtl_pc = spc65_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(65*4)]   <= 1'b0;
                  active_thread[(65*4)+1] <= 1'b0;
                  active_thread[(65*4)+2] <= 1'b0;
                  active_thread[(65*4)+3] <= 1'b0;
                  spc65_inst_done         <= 0;
                  spc65_phy_pc_w          <= 0;
                end else begin
                  active_thread[(65*4)]   <= 1'b1;
                  active_thread[(65*4)+1] <= 1'b1;
                  active_thread[(65*4)+2] <= 1'b1;
                  active_thread[(65*4)+3] <= 1'b1;
                  spc65_inst_done         <= `TILE65.piton_pc_vld;
                  spc65_phy_pc_w          <= `TILE65.piton_pc;
                end
            end
    

            assign spc66_thread_id = 2'b00;
            assign spc66_rtl_pc = spc66_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(66*4)]   <= 1'b0;
                  active_thread[(66*4)+1] <= 1'b0;
                  active_thread[(66*4)+2] <= 1'b0;
                  active_thread[(66*4)+3] <= 1'b0;
                  spc66_inst_done         <= 0;
                  spc66_phy_pc_w          <= 0;
                end else begin
                  active_thread[(66*4)]   <= 1'b1;
                  active_thread[(66*4)+1] <= 1'b1;
                  active_thread[(66*4)+2] <= 1'b1;
                  active_thread[(66*4)+3] <= 1'b1;
                  spc66_inst_done         <= `TILE66.piton_pc_vld;
                  spc66_phy_pc_w          <= `TILE66.piton_pc;
                end
            end
    

            assign spc67_thread_id = 2'b00;
            assign spc67_rtl_pc = spc67_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(67*4)]   <= 1'b0;
                  active_thread[(67*4)+1] <= 1'b0;
                  active_thread[(67*4)+2] <= 1'b0;
                  active_thread[(67*4)+3] <= 1'b0;
                  spc67_inst_done         <= 0;
                  spc67_phy_pc_w          <= 0;
                end else begin
                  active_thread[(67*4)]   <= 1'b1;
                  active_thread[(67*4)+1] <= 1'b1;
                  active_thread[(67*4)+2] <= 1'b1;
                  active_thread[(67*4)+3] <= 1'b1;
                  spc67_inst_done         <= `TILE67.piton_pc_vld;
                  spc67_phy_pc_w          <= `TILE67.piton_pc;
                end
            end
    

            assign spc68_thread_id = 2'b00;
            assign spc68_rtl_pc = spc68_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(68*4)]   <= 1'b0;
                  active_thread[(68*4)+1] <= 1'b0;
                  active_thread[(68*4)+2] <= 1'b0;
                  active_thread[(68*4)+3] <= 1'b0;
                  spc68_inst_done         <= 0;
                  spc68_phy_pc_w          <= 0;
                end else begin
                  active_thread[(68*4)]   <= 1'b1;
                  active_thread[(68*4)+1] <= 1'b1;
                  active_thread[(68*4)+2] <= 1'b1;
                  active_thread[(68*4)+3] <= 1'b1;
                  spc68_inst_done         <= `TILE68.piton_pc_vld;
                  spc68_phy_pc_w          <= `TILE68.piton_pc;
                end
            end
    

            assign spc69_thread_id = 2'b00;
            assign spc69_rtl_pc = spc69_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(69*4)]   <= 1'b0;
                  active_thread[(69*4)+1] <= 1'b0;
                  active_thread[(69*4)+2] <= 1'b0;
                  active_thread[(69*4)+3] <= 1'b0;
                  spc69_inst_done         <= 0;
                  spc69_phy_pc_w          <= 0;
                end else begin
                  active_thread[(69*4)]   <= 1'b1;
                  active_thread[(69*4)+1] <= 1'b1;
                  active_thread[(69*4)+2] <= 1'b1;
                  active_thread[(69*4)+3] <= 1'b1;
                  spc69_inst_done         <= `TILE69.piton_pc_vld;
                  spc69_phy_pc_w          <= `TILE69.piton_pc;
                end
            end
    

            assign spc70_thread_id = 2'b00;
            assign spc70_rtl_pc = spc70_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(70*4)]   <= 1'b0;
                  active_thread[(70*4)+1] <= 1'b0;
                  active_thread[(70*4)+2] <= 1'b0;
                  active_thread[(70*4)+3] <= 1'b0;
                  spc70_inst_done         <= 0;
                  spc70_phy_pc_w          <= 0;
                end else begin
                  active_thread[(70*4)]   <= 1'b1;
                  active_thread[(70*4)+1] <= 1'b1;
                  active_thread[(70*4)+2] <= 1'b1;
                  active_thread[(70*4)+3] <= 1'b1;
                  spc70_inst_done         <= `TILE70.piton_pc_vld;
                  spc70_phy_pc_w          <= `TILE70.piton_pc;
                end
            end
    

            assign spc71_thread_id = 2'b00;
            assign spc71_rtl_pc = spc71_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(71*4)]   <= 1'b0;
                  active_thread[(71*4)+1] <= 1'b0;
                  active_thread[(71*4)+2] <= 1'b0;
                  active_thread[(71*4)+3] <= 1'b0;
                  spc71_inst_done         <= 0;
                  spc71_phy_pc_w          <= 0;
                end else begin
                  active_thread[(71*4)]   <= 1'b1;
                  active_thread[(71*4)+1] <= 1'b1;
                  active_thread[(71*4)+2] <= 1'b1;
                  active_thread[(71*4)+3] <= 1'b1;
                  spc71_inst_done         <= `TILE71.piton_pc_vld;
                  spc71_phy_pc_w          <= `TILE71.piton_pc;
                end
            end
    

            assign spc72_thread_id = 2'b00;
            assign spc72_rtl_pc = spc72_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(72*4)]   <= 1'b0;
                  active_thread[(72*4)+1] <= 1'b0;
                  active_thread[(72*4)+2] <= 1'b0;
                  active_thread[(72*4)+3] <= 1'b0;
                  spc72_inst_done         <= 0;
                  spc72_phy_pc_w          <= 0;
                end else begin
                  active_thread[(72*4)]   <= 1'b1;
                  active_thread[(72*4)+1] <= 1'b1;
                  active_thread[(72*4)+2] <= 1'b1;
                  active_thread[(72*4)+3] <= 1'b1;
                  spc72_inst_done         <= `TILE72.piton_pc_vld;
                  spc72_phy_pc_w          <= `TILE72.piton_pc;
                end
            end
    

            assign spc73_thread_id = 2'b00;
            assign spc73_rtl_pc = spc73_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(73*4)]   <= 1'b0;
                  active_thread[(73*4)+1] <= 1'b0;
                  active_thread[(73*4)+2] <= 1'b0;
                  active_thread[(73*4)+3] <= 1'b0;
                  spc73_inst_done         <= 0;
                  spc73_phy_pc_w          <= 0;
                end else begin
                  active_thread[(73*4)]   <= 1'b1;
                  active_thread[(73*4)+1] <= 1'b1;
                  active_thread[(73*4)+2] <= 1'b1;
                  active_thread[(73*4)+3] <= 1'b1;
                  spc73_inst_done         <= `TILE73.piton_pc_vld;
                  spc73_phy_pc_w          <= `TILE73.piton_pc;
                end
            end
    

            assign spc74_thread_id = 2'b00;
            assign spc74_rtl_pc = spc74_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(74*4)]   <= 1'b0;
                  active_thread[(74*4)+1] <= 1'b0;
                  active_thread[(74*4)+2] <= 1'b0;
                  active_thread[(74*4)+3] <= 1'b0;
                  spc74_inst_done         <= 0;
                  spc74_phy_pc_w          <= 0;
                end else begin
                  active_thread[(74*4)]   <= 1'b1;
                  active_thread[(74*4)+1] <= 1'b1;
                  active_thread[(74*4)+2] <= 1'b1;
                  active_thread[(74*4)+3] <= 1'b1;
                  spc74_inst_done         <= `TILE74.piton_pc_vld;
                  spc74_phy_pc_w          <= `TILE74.piton_pc;
                end
            end
    

            assign spc75_thread_id = 2'b00;
            assign spc75_rtl_pc = spc75_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(75*4)]   <= 1'b0;
                  active_thread[(75*4)+1] <= 1'b0;
                  active_thread[(75*4)+2] <= 1'b0;
                  active_thread[(75*4)+3] <= 1'b0;
                  spc75_inst_done         <= 0;
                  spc75_phy_pc_w          <= 0;
                end else begin
                  active_thread[(75*4)]   <= 1'b1;
                  active_thread[(75*4)+1] <= 1'b1;
                  active_thread[(75*4)+2] <= 1'b1;
                  active_thread[(75*4)+3] <= 1'b1;
                  spc75_inst_done         <= `TILE75.piton_pc_vld;
                  spc75_phy_pc_w          <= `TILE75.piton_pc;
                end
            end
    

            assign spc76_thread_id = 2'b00;
            assign spc76_rtl_pc = spc76_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(76*4)]   <= 1'b0;
                  active_thread[(76*4)+1] <= 1'b0;
                  active_thread[(76*4)+2] <= 1'b0;
                  active_thread[(76*4)+3] <= 1'b0;
                  spc76_inst_done         <= 0;
                  spc76_phy_pc_w          <= 0;
                end else begin
                  active_thread[(76*4)]   <= 1'b1;
                  active_thread[(76*4)+1] <= 1'b1;
                  active_thread[(76*4)+2] <= 1'b1;
                  active_thread[(76*4)+3] <= 1'b1;
                  spc76_inst_done         <= `TILE76.piton_pc_vld;
                  spc76_phy_pc_w          <= `TILE76.piton_pc;
                end
            end
    

            assign spc77_thread_id = 2'b00;
            assign spc77_rtl_pc = spc77_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(77*4)]   <= 1'b0;
                  active_thread[(77*4)+1] <= 1'b0;
                  active_thread[(77*4)+2] <= 1'b0;
                  active_thread[(77*4)+3] <= 1'b0;
                  spc77_inst_done         <= 0;
                  spc77_phy_pc_w          <= 0;
                end else begin
                  active_thread[(77*4)]   <= 1'b1;
                  active_thread[(77*4)+1] <= 1'b1;
                  active_thread[(77*4)+2] <= 1'b1;
                  active_thread[(77*4)+3] <= 1'b1;
                  spc77_inst_done         <= `TILE77.piton_pc_vld;
                  spc77_phy_pc_w          <= `TILE77.piton_pc;
                end
            end
    

            assign spc78_thread_id = 2'b00;
            assign spc78_rtl_pc = spc78_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(78*4)]   <= 1'b0;
                  active_thread[(78*4)+1] <= 1'b0;
                  active_thread[(78*4)+2] <= 1'b0;
                  active_thread[(78*4)+3] <= 1'b0;
                  spc78_inst_done         <= 0;
                  spc78_phy_pc_w          <= 0;
                end else begin
                  active_thread[(78*4)]   <= 1'b1;
                  active_thread[(78*4)+1] <= 1'b1;
                  active_thread[(78*4)+2] <= 1'b1;
                  active_thread[(78*4)+3] <= 1'b1;
                  spc78_inst_done         <= `TILE78.piton_pc_vld;
                  spc78_phy_pc_w          <= `TILE78.piton_pc;
                end
            end
    

            assign spc79_thread_id = 2'b00;
            assign spc79_rtl_pc = spc79_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(79*4)]   <= 1'b0;
                  active_thread[(79*4)+1] <= 1'b0;
                  active_thread[(79*4)+2] <= 1'b0;
                  active_thread[(79*4)+3] <= 1'b0;
                  spc79_inst_done         <= 0;
                  spc79_phy_pc_w          <= 0;
                end else begin
                  active_thread[(79*4)]   <= 1'b1;
                  active_thread[(79*4)+1] <= 1'b1;
                  active_thread[(79*4)+2] <= 1'b1;
                  active_thread[(79*4)+3] <= 1'b1;
                  spc79_inst_done         <= `TILE79.piton_pc_vld;
                  spc79_phy_pc_w          <= `TILE79.piton_pc;
                end
            end
    

            assign spc80_thread_id = 2'b00;
            assign spc80_rtl_pc = spc80_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(80*4)]   <= 1'b0;
                  active_thread[(80*4)+1] <= 1'b0;
                  active_thread[(80*4)+2] <= 1'b0;
                  active_thread[(80*4)+3] <= 1'b0;
                  spc80_inst_done         <= 0;
                  spc80_phy_pc_w          <= 0;
                end else begin
                  active_thread[(80*4)]   <= 1'b1;
                  active_thread[(80*4)+1] <= 1'b1;
                  active_thread[(80*4)+2] <= 1'b1;
                  active_thread[(80*4)+3] <= 1'b1;
                  spc80_inst_done         <= `TILE80.piton_pc_vld;
                  spc80_phy_pc_w          <= `TILE80.piton_pc;
                end
            end
    

            assign spc81_thread_id = 2'b00;
            assign spc81_rtl_pc = spc81_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(81*4)]   <= 1'b0;
                  active_thread[(81*4)+1] <= 1'b0;
                  active_thread[(81*4)+2] <= 1'b0;
                  active_thread[(81*4)+3] <= 1'b0;
                  spc81_inst_done         <= 0;
                  spc81_phy_pc_w          <= 0;
                end else begin
                  active_thread[(81*4)]   <= 1'b1;
                  active_thread[(81*4)+1] <= 1'b1;
                  active_thread[(81*4)+2] <= 1'b1;
                  active_thread[(81*4)+3] <= 1'b1;
                  spc81_inst_done         <= `TILE81.piton_pc_vld;
                  spc81_phy_pc_w          <= `TILE81.piton_pc;
                end
            end
    

            assign spc82_thread_id = 2'b00;
            assign spc82_rtl_pc = spc82_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(82*4)]   <= 1'b0;
                  active_thread[(82*4)+1] <= 1'b0;
                  active_thread[(82*4)+2] <= 1'b0;
                  active_thread[(82*4)+3] <= 1'b0;
                  spc82_inst_done         <= 0;
                  spc82_phy_pc_w          <= 0;
                end else begin
                  active_thread[(82*4)]   <= 1'b1;
                  active_thread[(82*4)+1] <= 1'b1;
                  active_thread[(82*4)+2] <= 1'b1;
                  active_thread[(82*4)+3] <= 1'b1;
                  spc82_inst_done         <= `TILE82.piton_pc_vld;
                  spc82_phy_pc_w          <= `TILE82.piton_pc;
                end
            end
    

            assign spc83_thread_id = 2'b00;
            assign spc83_rtl_pc = spc83_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(83*4)]   <= 1'b0;
                  active_thread[(83*4)+1] <= 1'b0;
                  active_thread[(83*4)+2] <= 1'b0;
                  active_thread[(83*4)+3] <= 1'b0;
                  spc83_inst_done         <= 0;
                  spc83_phy_pc_w          <= 0;
                end else begin
                  active_thread[(83*4)]   <= 1'b1;
                  active_thread[(83*4)+1] <= 1'b1;
                  active_thread[(83*4)+2] <= 1'b1;
                  active_thread[(83*4)+3] <= 1'b1;
                  spc83_inst_done         <= `TILE83.piton_pc_vld;
                  spc83_phy_pc_w          <= `TILE83.piton_pc;
                end
            end
    

            assign spc84_thread_id = 2'b00;
            assign spc84_rtl_pc = spc84_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(84*4)]   <= 1'b0;
                  active_thread[(84*4)+1] <= 1'b0;
                  active_thread[(84*4)+2] <= 1'b0;
                  active_thread[(84*4)+3] <= 1'b0;
                  spc84_inst_done         <= 0;
                  spc84_phy_pc_w          <= 0;
                end else begin
                  active_thread[(84*4)]   <= 1'b1;
                  active_thread[(84*4)+1] <= 1'b1;
                  active_thread[(84*4)+2] <= 1'b1;
                  active_thread[(84*4)+3] <= 1'b1;
                  spc84_inst_done         <= `TILE84.piton_pc_vld;
                  spc84_phy_pc_w          <= `TILE84.piton_pc;
                end
            end
    

            assign spc85_thread_id = 2'b00;
            assign spc85_rtl_pc = spc85_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(85*4)]   <= 1'b0;
                  active_thread[(85*4)+1] <= 1'b0;
                  active_thread[(85*4)+2] <= 1'b0;
                  active_thread[(85*4)+3] <= 1'b0;
                  spc85_inst_done         <= 0;
                  spc85_phy_pc_w          <= 0;
                end else begin
                  active_thread[(85*4)]   <= 1'b1;
                  active_thread[(85*4)+1] <= 1'b1;
                  active_thread[(85*4)+2] <= 1'b1;
                  active_thread[(85*4)+3] <= 1'b1;
                  spc85_inst_done         <= `TILE85.piton_pc_vld;
                  spc85_phy_pc_w          <= `TILE85.piton_pc;
                end
            end
    

            assign spc86_thread_id = 2'b00;
            assign spc86_rtl_pc = spc86_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(86*4)]   <= 1'b0;
                  active_thread[(86*4)+1] <= 1'b0;
                  active_thread[(86*4)+2] <= 1'b0;
                  active_thread[(86*4)+3] <= 1'b0;
                  spc86_inst_done         <= 0;
                  spc86_phy_pc_w          <= 0;
                end else begin
                  active_thread[(86*4)]   <= 1'b1;
                  active_thread[(86*4)+1] <= 1'b1;
                  active_thread[(86*4)+2] <= 1'b1;
                  active_thread[(86*4)+3] <= 1'b1;
                  spc86_inst_done         <= `TILE86.piton_pc_vld;
                  spc86_phy_pc_w          <= `TILE86.piton_pc;
                end
            end
    

            assign spc87_thread_id = 2'b00;
            assign spc87_rtl_pc = spc87_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(87*4)]   <= 1'b0;
                  active_thread[(87*4)+1] <= 1'b0;
                  active_thread[(87*4)+2] <= 1'b0;
                  active_thread[(87*4)+3] <= 1'b0;
                  spc87_inst_done         <= 0;
                  spc87_phy_pc_w          <= 0;
                end else begin
                  active_thread[(87*4)]   <= 1'b1;
                  active_thread[(87*4)+1] <= 1'b1;
                  active_thread[(87*4)+2] <= 1'b1;
                  active_thread[(87*4)+3] <= 1'b1;
                  spc87_inst_done         <= `TILE87.piton_pc_vld;
                  spc87_phy_pc_w          <= `TILE87.piton_pc;
                end
            end
    

            assign spc88_thread_id = 2'b00;
            assign spc88_rtl_pc = spc88_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(88*4)]   <= 1'b0;
                  active_thread[(88*4)+1] <= 1'b0;
                  active_thread[(88*4)+2] <= 1'b0;
                  active_thread[(88*4)+3] <= 1'b0;
                  spc88_inst_done         <= 0;
                  spc88_phy_pc_w          <= 0;
                end else begin
                  active_thread[(88*4)]   <= 1'b1;
                  active_thread[(88*4)+1] <= 1'b1;
                  active_thread[(88*4)+2] <= 1'b1;
                  active_thread[(88*4)+3] <= 1'b1;
                  spc88_inst_done         <= `TILE88.piton_pc_vld;
                  spc88_phy_pc_w          <= `TILE88.piton_pc;
                end
            end
    

            assign spc89_thread_id = 2'b00;
            assign spc89_rtl_pc = spc89_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(89*4)]   <= 1'b0;
                  active_thread[(89*4)+1] <= 1'b0;
                  active_thread[(89*4)+2] <= 1'b0;
                  active_thread[(89*4)+3] <= 1'b0;
                  spc89_inst_done         <= 0;
                  spc89_phy_pc_w          <= 0;
                end else begin
                  active_thread[(89*4)]   <= 1'b1;
                  active_thread[(89*4)+1] <= 1'b1;
                  active_thread[(89*4)+2] <= 1'b1;
                  active_thread[(89*4)+3] <= 1'b1;
                  spc89_inst_done         <= `TILE89.piton_pc_vld;
                  spc89_phy_pc_w          <= `TILE89.piton_pc;
                end
            end
    

            assign spc90_thread_id = 2'b00;
            assign spc90_rtl_pc = spc90_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(90*4)]   <= 1'b0;
                  active_thread[(90*4)+1] <= 1'b0;
                  active_thread[(90*4)+2] <= 1'b0;
                  active_thread[(90*4)+3] <= 1'b0;
                  spc90_inst_done         <= 0;
                  spc90_phy_pc_w          <= 0;
                end else begin
                  active_thread[(90*4)]   <= 1'b1;
                  active_thread[(90*4)+1] <= 1'b1;
                  active_thread[(90*4)+2] <= 1'b1;
                  active_thread[(90*4)+3] <= 1'b1;
                  spc90_inst_done         <= `TILE90.piton_pc_vld;
                  spc90_phy_pc_w          <= `TILE90.piton_pc;
                end
            end
    

            assign spc91_thread_id = 2'b00;
            assign spc91_rtl_pc = spc91_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(91*4)]   <= 1'b0;
                  active_thread[(91*4)+1] <= 1'b0;
                  active_thread[(91*4)+2] <= 1'b0;
                  active_thread[(91*4)+3] <= 1'b0;
                  spc91_inst_done         <= 0;
                  spc91_phy_pc_w          <= 0;
                end else begin
                  active_thread[(91*4)]   <= 1'b1;
                  active_thread[(91*4)+1] <= 1'b1;
                  active_thread[(91*4)+2] <= 1'b1;
                  active_thread[(91*4)+3] <= 1'b1;
                  spc91_inst_done         <= `TILE91.piton_pc_vld;
                  spc91_phy_pc_w          <= `TILE91.piton_pc;
                end
            end
    

            assign spc92_thread_id = 2'b00;
            assign spc92_rtl_pc = spc92_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(92*4)]   <= 1'b0;
                  active_thread[(92*4)+1] <= 1'b0;
                  active_thread[(92*4)+2] <= 1'b0;
                  active_thread[(92*4)+3] <= 1'b0;
                  spc92_inst_done         <= 0;
                  spc92_phy_pc_w          <= 0;
                end else begin
                  active_thread[(92*4)]   <= 1'b1;
                  active_thread[(92*4)+1] <= 1'b1;
                  active_thread[(92*4)+2] <= 1'b1;
                  active_thread[(92*4)+3] <= 1'b1;
                  spc92_inst_done         <= `TILE92.piton_pc_vld;
                  spc92_phy_pc_w          <= `TILE92.piton_pc;
                end
            end
    

            assign spc93_thread_id = 2'b00;
            assign spc93_rtl_pc = spc93_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(93*4)]   <= 1'b0;
                  active_thread[(93*4)+1] <= 1'b0;
                  active_thread[(93*4)+2] <= 1'b0;
                  active_thread[(93*4)+3] <= 1'b0;
                  spc93_inst_done         <= 0;
                  spc93_phy_pc_w          <= 0;
                end else begin
                  active_thread[(93*4)]   <= 1'b1;
                  active_thread[(93*4)+1] <= 1'b1;
                  active_thread[(93*4)+2] <= 1'b1;
                  active_thread[(93*4)+3] <= 1'b1;
                  spc93_inst_done         <= `TILE93.piton_pc_vld;
                  spc93_phy_pc_w          <= `TILE93.piton_pc;
                end
            end
    

            assign spc94_thread_id = 2'b00;
            assign spc94_rtl_pc = spc94_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(94*4)]   <= 1'b0;
                  active_thread[(94*4)+1] <= 1'b0;
                  active_thread[(94*4)+2] <= 1'b0;
                  active_thread[(94*4)+3] <= 1'b0;
                  spc94_inst_done         <= 0;
                  spc94_phy_pc_w          <= 0;
                end else begin
                  active_thread[(94*4)]   <= 1'b1;
                  active_thread[(94*4)+1] <= 1'b1;
                  active_thread[(94*4)+2] <= 1'b1;
                  active_thread[(94*4)+3] <= 1'b1;
                  spc94_inst_done         <= `TILE94.piton_pc_vld;
                  spc94_phy_pc_w          <= `TILE94.piton_pc;
                end
            end
    

            assign spc95_thread_id = 2'b00;
            assign spc95_rtl_pc = spc95_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(95*4)]   <= 1'b0;
                  active_thread[(95*4)+1] <= 1'b0;
                  active_thread[(95*4)+2] <= 1'b0;
                  active_thread[(95*4)+3] <= 1'b0;
                  spc95_inst_done         <= 0;
                  spc95_phy_pc_w          <= 0;
                end else begin
                  active_thread[(95*4)]   <= 1'b1;
                  active_thread[(95*4)+1] <= 1'b1;
                  active_thread[(95*4)+2] <= 1'b1;
                  active_thread[(95*4)+3] <= 1'b1;
                  spc95_inst_done         <= `TILE95.piton_pc_vld;
                  spc95_phy_pc_w          <= `TILE95.piton_pc;
                end
            end
    

            assign spc96_thread_id = 2'b00;
            assign spc96_rtl_pc = spc96_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(96*4)]   <= 1'b0;
                  active_thread[(96*4)+1] <= 1'b0;
                  active_thread[(96*4)+2] <= 1'b0;
                  active_thread[(96*4)+3] <= 1'b0;
                  spc96_inst_done         <= 0;
                  spc96_phy_pc_w          <= 0;
                end else begin
                  active_thread[(96*4)]   <= 1'b1;
                  active_thread[(96*4)+1] <= 1'b1;
                  active_thread[(96*4)+2] <= 1'b1;
                  active_thread[(96*4)+3] <= 1'b1;
                  spc96_inst_done         <= `TILE96.piton_pc_vld;
                  spc96_phy_pc_w          <= `TILE96.piton_pc;
                end
            end
    

            assign spc97_thread_id = 2'b00;
            assign spc97_rtl_pc = spc97_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(97*4)]   <= 1'b0;
                  active_thread[(97*4)+1] <= 1'b0;
                  active_thread[(97*4)+2] <= 1'b0;
                  active_thread[(97*4)+3] <= 1'b0;
                  spc97_inst_done         <= 0;
                  spc97_phy_pc_w          <= 0;
                end else begin
                  active_thread[(97*4)]   <= 1'b1;
                  active_thread[(97*4)+1] <= 1'b1;
                  active_thread[(97*4)+2] <= 1'b1;
                  active_thread[(97*4)+3] <= 1'b1;
                  spc97_inst_done         <= `TILE97.piton_pc_vld;
                  spc97_phy_pc_w          <= `TILE97.piton_pc;
                end
            end
    

            assign spc98_thread_id = 2'b00;
            assign spc98_rtl_pc = spc98_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(98*4)]   <= 1'b0;
                  active_thread[(98*4)+1] <= 1'b0;
                  active_thread[(98*4)+2] <= 1'b0;
                  active_thread[(98*4)+3] <= 1'b0;
                  spc98_inst_done         <= 0;
                  spc98_phy_pc_w          <= 0;
                end else begin
                  active_thread[(98*4)]   <= 1'b1;
                  active_thread[(98*4)+1] <= 1'b1;
                  active_thread[(98*4)+2] <= 1'b1;
                  active_thread[(98*4)+3] <= 1'b1;
                  spc98_inst_done         <= `TILE98.piton_pc_vld;
                  spc98_phy_pc_w          <= `TILE98.piton_pc;
                end
            end
    

            assign spc99_thread_id = 2'b00;
            assign spc99_rtl_pc = spc99_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(99*4)]   <= 1'b0;
                  active_thread[(99*4)+1] <= 1'b0;
                  active_thread[(99*4)+2] <= 1'b0;
                  active_thread[(99*4)+3] <= 1'b0;
                  spc99_inst_done         <= 0;
                  spc99_phy_pc_w          <= 0;
                end else begin
                  active_thread[(99*4)]   <= 1'b1;
                  active_thread[(99*4)+1] <= 1'b1;
                  active_thread[(99*4)+2] <= 1'b1;
                  active_thread[(99*4)+3] <= 1'b1;
                  spc99_inst_done         <= `TILE99.piton_pc_vld;
                  spc99_phy_pc_w          <= `TILE99.piton_pc;
                end
            end
    

            assign spc100_thread_id = 2'b00;
            assign spc100_rtl_pc = spc100_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(100*4)]   <= 1'b0;
                  active_thread[(100*4)+1] <= 1'b0;
                  active_thread[(100*4)+2] <= 1'b0;
                  active_thread[(100*4)+3] <= 1'b0;
                  spc100_inst_done         <= 0;
                  spc100_phy_pc_w          <= 0;
                end else begin
                  active_thread[(100*4)]   <= 1'b1;
                  active_thread[(100*4)+1] <= 1'b1;
                  active_thread[(100*4)+2] <= 1'b1;
                  active_thread[(100*4)+3] <= 1'b1;
                  spc100_inst_done         <= `TILE100.piton_pc_vld;
                  spc100_phy_pc_w          <= `TILE100.piton_pc;
                end
            end
    

            assign spc101_thread_id = 2'b00;
            assign spc101_rtl_pc = spc101_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(101*4)]   <= 1'b0;
                  active_thread[(101*4)+1] <= 1'b0;
                  active_thread[(101*4)+2] <= 1'b0;
                  active_thread[(101*4)+3] <= 1'b0;
                  spc101_inst_done         <= 0;
                  spc101_phy_pc_w          <= 0;
                end else begin
                  active_thread[(101*4)]   <= 1'b1;
                  active_thread[(101*4)+1] <= 1'b1;
                  active_thread[(101*4)+2] <= 1'b1;
                  active_thread[(101*4)+3] <= 1'b1;
                  spc101_inst_done         <= `TILE101.piton_pc_vld;
                  spc101_phy_pc_w          <= `TILE101.piton_pc;
                end
            end
    

            assign spc102_thread_id = 2'b00;
            assign spc102_rtl_pc = spc102_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(102*4)]   <= 1'b0;
                  active_thread[(102*4)+1] <= 1'b0;
                  active_thread[(102*4)+2] <= 1'b0;
                  active_thread[(102*4)+3] <= 1'b0;
                  spc102_inst_done         <= 0;
                  spc102_phy_pc_w          <= 0;
                end else begin
                  active_thread[(102*4)]   <= 1'b1;
                  active_thread[(102*4)+1] <= 1'b1;
                  active_thread[(102*4)+2] <= 1'b1;
                  active_thread[(102*4)+3] <= 1'b1;
                  spc102_inst_done         <= `TILE102.piton_pc_vld;
                  spc102_phy_pc_w          <= `TILE102.piton_pc;
                end
            end
    

            assign spc103_thread_id = 2'b00;
            assign spc103_rtl_pc = spc103_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(103*4)]   <= 1'b0;
                  active_thread[(103*4)+1] <= 1'b0;
                  active_thread[(103*4)+2] <= 1'b0;
                  active_thread[(103*4)+3] <= 1'b0;
                  spc103_inst_done         <= 0;
                  spc103_phy_pc_w          <= 0;
                end else begin
                  active_thread[(103*4)]   <= 1'b1;
                  active_thread[(103*4)+1] <= 1'b1;
                  active_thread[(103*4)+2] <= 1'b1;
                  active_thread[(103*4)+3] <= 1'b1;
                  spc103_inst_done         <= `TILE103.piton_pc_vld;
                  spc103_phy_pc_w          <= `TILE103.piton_pc;
                end
            end
    

            assign spc104_thread_id = 2'b00;
            assign spc104_rtl_pc = spc104_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(104*4)]   <= 1'b0;
                  active_thread[(104*4)+1] <= 1'b0;
                  active_thread[(104*4)+2] <= 1'b0;
                  active_thread[(104*4)+3] <= 1'b0;
                  spc104_inst_done         <= 0;
                  spc104_phy_pc_w          <= 0;
                end else begin
                  active_thread[(104*4)]   <= 1'b1;
                  active_thread[(104*4)+1] <= 1'b1;
                  active_thread[(104*4)+2] <= 1'b1;
                  active_thread[(104*4)+3] <= 1'b1;
                  spc104_inst_done         <= `TILE104.piton_pc_vld;
                  spc104_phy_pc_w          <= `TILE104.piton_pc;
                end
            end
    

            assign spc105_thread_id = 2'b00;
            assign spc105_rtl_pc = spc105_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(105*4)]   <= 1'b0;
                  active_thread[(105*4)+1] <= 1'b0;
                  active_thread[(105*4)+2] <= 1'b0;
                  active_thread[(105*4)+3] <= 1'b0;
                  spc105_inst_done         <= 0;
                  spc105_phy_pc_w          <= 0;
                end else begin
                  active_thread[(105*4)]   <= 1'b1;
                  active_thread[(105*4)+1] <= 1'b1;
                  active_thread[(105*4)+2] <= 1'b1;
                  active_thread[(105*4)+3] <= 1'b1;
                  spc105_inst_done         <= `TILE105.piton_pc_vld;
                  spc105_phy_pc_w          <= `TILE105.piton_pc;
                end
            end
    

            assign spc106_thread_id = 2'b00;
            assign spc106_rtl_pc = spc106_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(106*4)]   <= 1'b0;
                  active_thread[(106*4)+1] <= 1'b0;
                  active_thread[(106*4)+2] <= 1'b0;
                  active_thread[(106*4)+3] <= 1'b0;
                  spc106_inst_done         <= 0;
                  spc106_phy_pc_w          <= 0;
                end else begin
                  active_thread[(106*4)]   <= 1'b1;
                  active_thread[(106*4)+1] <= 1'b1;
                  active_thread[(106*4)+2] <= 1'b1;
                  active_thread[(106*4)+3] <= 1'b1;
                  spc106_inst_done         <= `TILE106.piton_pc_vld;
                  spc106_phy_pc_w          <= `TILE106.piton_pc;
                end
            end
    

            assign spc107_thread_id = 2'b00;
            assign spc107_rtl_pc = spc107_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(107*4)]   <= 1'b0;
                  active_thread[(107*4)+1] <= 1'b0;
                  active_thread[(107*4)+2] <= 1'b0;
                  active_thread[(107*4)+3] <= 1'b0;
                  spc107_inst_done         <= 0;
                  spc107_phy_pc_w          <= 0;
                end else begin
                  active_thread[(107*4)]   <= 1'b1;
                  active_thread[(107*4)+1] <= 1'b1;
                  active_thread[(107*4)+2] <= 1'b1;
                  active_thread[(107*4)+3] <= 1'b1;
                  spc107_inst_done         <= `TILE107.piton_pc_vld;
                  spc107_phy_pc_w          <= `TILE107.piton_pc;
                end
            end
    

            assign spc108_thread_id = 2'b00;
            assign spc108_rtl_pc = spc108_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(108*4)]   <= 1'b0;
                  active_thread[(108*4)+1] <= 1'b0;
                  active_thread[(108*4)+2] <= 1'b0;
                  active_thread[(108*4)+3] <= 1'b0;
                  spc108_inst_done         <= 0;
                  spc108_phy_pc_w          <= 0;
                end else begin
                  active_thread[(108*4)]   <= 1'b1;
                  active_thread[(108*4)+1] <= 1'b1;
                  active_thread[(108*4)+2] <= 1'b1;
                  active_thread[(108*4)+3] <= 1'b1;
                  spc108_inst_done         <= `TILE108.piton_pc_vld;
                  spc108_phy_pc_w          <= `TILE108.piton_pc;
                end
            end
    

            assign spc109_thread_id = 2'b00;
            assign spc109_rtl_pc = spc109_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(109*4)]   <= 1'b0;
                  active_thread[(109*4)+1] <= 1'b0;
                  active_thread[(109*4)+2] <= 1'b0;
                  active_thread[(109*4)+3] <= 1'b0;
                  spc109_inst_done         <= 0;
                  spc109_phy_pc_w          <= 0;
                end else begin
                  active_thread[(109*4)]   <= 1'b1;
                  active_thread[(109*4)+1] <= 1'b1;
                  active_thread[(109*4)+2] <= 1'b1;
                  active_thread[(109*4)+3] <= 1'b1;
                  spc109_inst_done         <= `TILE109.piton_pc_vld;
                  spc109_phy_pc_w          <= `TILE109.piton_pc;
                end
            end
    

            assign spc110_thread_id = 2'b00;
            assign spc110_rtl_pc = spc110_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(110*4)]   <= 1'b0;
                  active_thread[(110*4)+1] <= 1'b0;
                  active_thread[(110*4)+2] <= 1'b0;
                  active_thread[(110*4)+3] <= 1'b0;
                  spc110_inst_done         <= 0;
                  spc110_phy_pc_w          <= 0;
                end else begin
                  active_thread[(110*4)]   <= 1'b1;
                  active_thread[(110*4)+1] <= 1'b1;
                  active_thread[(110*4)+2] <= 1'b1;
                  active_thread[(110*4)+3] <= 1'b1;
                  spc110_inst_done         <= `TILE110.piton_pc_vld;
                  spc110_phy_pc_w          <= `TILE110.piton_pc;
                end
            end
    

            assign spc111_thread_id = 2'b00;
            assign spc111_rtl_pc = spc111_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(111*4)]   <= 1'b0;
                  active_thread[(111*4)+1] <= 1'b0;
                  active_thread[(111*4)+2] <= 1'b0;
                  active_thread[(111*4)+3] <= 1'b0;
                  spc111_inst_done         <= 0;
                  spc111_phy_pc_w          <= 0;
                end else begin
                  active_thread[(111*4)]   <= 1'b1;
                  active_thread[(111*4)+1] <= 1'b1;
                  active_thread[(111*4)+2] <= 1'b1;
                  active_thread[(111*4)+3] <= 1'b1;
                  spc111_inst_done         <= `TILE111.piton_pc_vld;
                  spc111_phy_pc_w          <= `TILE111.piton_pc;
                end
            end
    

            assign spc112_thread_id = 2'b00;
            assign spc112_rtl_pc = spc112_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(112*4)]   <= 1'b0;
                  active_thread[(112*4)+1] <= 1'b0;
                  active_thread[(112*4)+2] <= 1'b0;
                  active_thread[(112*4)+3] <= 1'b0;
                  spc112_inst_done         <= 0;
                  spc112_phy_pc_w          <= 0;
                end else begin
                  active_thread[(112*4)]   <= 1'b1;
                  active_thread[(112*4)+1] <= 1'b1;
                  active_thread[(112*4)+2] <= 1'b1;
                  active_thread[(112*4)+3] <= 1'b1;
                  spc112_inst_done         <= `TILE112.piton_pc_vld;
                  spc112_phy_pc_w          <= `TILE112.piton_pc;
                end
            end
    

            assign spc113_thread_id = 2'b00;
            assign spc113_rtl_pc = spc113_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(113*4)]   <= 1'b0;
                  active_thread[(113*4)+1] <= 1'b0;
                  active_thread[(113*4)+2] <= 1'b0;
                  active_thread[(113*4)+3] <= 1'b0;
                  spc113_inst_done         <= 0;
                  spc113_phy_pc_w          <= 0;
                end else begin
                  active_thread[(113*4)]   <= 1'b1;
                  active_thread[(113*4)+1] <= 1'b1;
                  active_thread[(113*4)+2] <= 1'b1;
                  active_thread[(113*4)+3] <= 1'b1;
                  spc113_inst_done         <= `TILE113.piton_pc_vld;
                  spc113_phy_pc_w          <= `TILE113.piton_pc;
                end
            end
    

            assign spc114_thread_id = 2'b00;
            assign spc114_rtl_pc = spc114_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(114*4)]   <= 1'b0;
                  active_thread[(114*4)+1] <= 1'b0;
                  active_thread[(114*4)+2] <= 1'b0;
                  active_thread[(114*4)+3] <= 1'b0;
                  spc114_inst_done         <= 0;
                  spc114_phy_pc_w          <= 0;
                end else begin
                  active_thread[(114*4)]   <= 1'b1;
                  active_thread[(114*4)+1] <= 1'b1;
                  active_thread[(114*4)+2] <= 1'b1;
                  active_thread[(114*4)+3] <= 1'b1;
                  spc114_inst_done         <= `TILE114.piton_pc_vld;
                  spc114_phy_pc_w          <= `TILE114.piton_pc;
                end
            end
    

            assign spc115_thread_id = 2'b00;
            assign spc115_rtl_pc = spc115_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(115*4)]   <= 1'b0;
                  active_thread[(115*4)+1] <= 1'b0;
                  active_thread[(115*4)+2] <= 1'b0;
                  active_thread[(115*4)+3] <= 1'b0;
                  spc115_inst_done         <= 0;
                  spc115_phy_pc_w          <= 0;
                end else begin
                  active_thread[(115*4)]   <= 1'b1;
                  active_thread[(115*4)+1] <= 1'b1;
                  active_thread[(115*4)+2] <= 1'b1;
                  active_thread[(115*4)+3] <= 1'b1;
                  spc115_inst_done         <= `TILE115.piton_pc_vld;
                  spc115_phy_pc_w          <= `TILE115.piton_pc;
                end
            end
    

            assign spc116_thread_id = 2'b00;
            assign spc116_rtl_pc = spc116_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(116*4)]   <= 1'b0;
                  active_thread[(116*4)+1] <= 1'b0;
                  active_thread[(116*4)+2] <= 1'b0;
                  active_thread[(116*4)+3] <= 1'b0;
                  spc116_inst_done         <= 0;
                  spc116_phy_pc_w          <= 0;
                end else begin
                  active_thread[(116*4)]   <= 1'b1;
                  active_thread[(116*4)+1] <= 1'b1;
                  active_thread[(116*4)+2] <= 1'b1;
                  active_thread[(116*4)+3] <= 1'b1;
                  spc116_inst_done         <= `TILE116.piton_pc_vld;
                  spc116_phy_pc_w          <= `TILE116.piton_pc;
                end
            end
    

            assign spc117_thread_id = 2'b00;
            assign spc117_rtl_pc = spc117_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(117*4)]   <= 1'b0;
                  active_thread[(117*4)+1] <= 1'b0;
                  active_thread[(117*4)+2] <= 1'b0;
                  active_thread[(117*4)+3] <= 1'b0;
                  spc117_inst_done         <= 0;
                  spc117_phy_pc_w          <= 0;
                end else begin
                  active_thread[(117*4)]   <= 1'b1;
                  active_thread[(117*4)+1] <= 1'b1;
                  active_thread[(117*4)+2] <= 1'b1;
                  active_thread[(117*4)+3] <= 1'b1;
                  spc117_inst_done         <= `TILE117.piton_pc_vld;
                  spc117_phy_pc_w          <= `TILE117.piton_pc;
                end
            end
    

            assign spc118_thread_id = 2'b00;
            assign spc118_rtl_pc = spc118_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(118*4)]   <= 1'b0;
                  active_thread[(118*4)+1] <= 1'b0;
                  active_thread[(118*4)+2] <= 1'b0;
                  active_thread[(118*4)+3] <= 1'b0;
                  spc118_inst_done         <= 0;
                  spc118_phy_pc_w          <= 0;
                end else begin
                  active_thread[(118*4)]   <= 1'b1;
                  active_thread[(118*4)+1] <= 1'b1;
                  active_thread[(118*4)+2] <= 1'b1;
                  active_thread[(118*4)+3] <= 1'b1;
                  spc118_inst_done         <= `TILE118.piton_pc_vld;
                  spc118_phy_pc_w          <= `TILE118.piton_pc;
                end
            end
    

            assign spc119_thread_id = 2'b00;
            assign spc119_rtl_pc = spc119_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(119*4)]   <= 1'b0;
                  active_thread[(119*4)+1] <= 1'b0;
                  active_thread[(119*4)+2] <= 1'b0;
                  active_thread[(119*4)+3] <= 1'b0;
                  spc119_inst_done         <= 0;
                  spc119_phy_pc_w          <= 0;
                end else begin
                  active_thread[(119*4)]   <= 1'b1;
                  active_thread[(119*4)+1] <= 1'b1;
                  active_thread[(119*4)+2] <= 1'b1;
                  active_thread[(119*4)+3] <= 1'b1;
                  spc119_inst_done         <= `TILE119.piton_pc_vld;
                  spc119_phy_pc_w          <= `TILE119.piton_pc;
                end
            end
    

            assign spc120_thread_id = 2'b00;
            assign spc120_rtl_pc = spc120_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(120*4)]   <= 1'b0;
                  active_thread[(120*4)+1] <= 1'b0;
                  active_thread[(120*4)+2] <= 1'b0;
                  active_thread[(120*4)+3] <= 1'b0;
                  spc120_inst_done         <= 0;
                  spc120_phy_pc_w          <= 0;
                end else begin
                  active_thread[(120*4)]   <= 1'b1;
                  active_thread[(120*4)+1] <= 1'b1;
                  active_thread[(120*4)+2] <= 1'b1;
                  active_thread[(120*4)+3] <= 1'b1;
                  spc120_inst_done         <= `TILE120.piton_pc_vld;
                  spc120_phy_pc_w          <= `TILE120.piton_pc;
                end
            end
    

            assign spc121_thread_id = 2'b00;
            assign spc121_rtl_pc = spc121_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(121*4)]   <= 1'b0;
                  active_thread[(121*4)+1] <= 1'b0;
                  active_thread[(121*4)+2] <= 1'b0;
                  active_thread[(121*4)+3] <= 1'b0;
                  spc121_inst_done         <= 0;
                  spc121_phy_pc_w          <= 0;
                end else begin
                  active_thread[(121*4)]   <= 1'b1;
                  active_thread[(121*4)+1] <= 1'b1;
                  active_thread[(121*4)+2] <= 1'b1;
                  active_thread[(121*4)+3] <= 1'b1;
                  spc121_inst_done         <= `TILE121.piton_pc_vld;
                  spc121_phy_pc_w          <= `TILE121.piton_pc;
                end
            end
    

            assign spc122_thread_id = 2'b00;
            assign spc122_rtl_pc = spc122_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(122*4)]   <= 1'b0;
                  active_thread[(122*4)+1] <= 1'b0;
                  active_thread[(122*4)+2] <= 1'b0;
                  active_thread[(122*4)+3] <= 1'b0;
                  spc122_inst_done         <= 0;
                  spc122_phy_pc_w          <= 0;
                end else begin
                  active_thread[(122*4)]   <= 1'b1;
                  active_thread[(122*4)+1] <= 1'b1;
                  active_thread[(122*4)+2] <= 1'b1;
                  active_thread[(122*4)+3] <= 1'b1;
                  spc122_inst_done         <= `TILE122.piton_pc_vld;
                  spc122_phy_pc_w          <= `TILE122.piton_pc;
                end
            end
    

            assign spc123_thread_id = 2'b00;
            assign spc123_rtl_pc = spc123_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(123*4)]   <= 1'b0;
                  active_thread[(123*4)+1] <= 1'b0;
                  active_thread[(123*4)+2] <= 1'b0;
                  active_thread[(123*4)+3] <= 1'b0;
                  spc123_inst_done         <= 0;
                  spc123_phy_pc_w          <= 0;
                end else begin
                  active_thread[(123*4)]   <= 1'b1;
                  active_thread[(123*4)+1] <= 1'b1;
                  active_thread[(123*4)+2] <= 1'b1;
                  active_thread[(123*4)+3] <= 1'b1;
                  spc123_inst_done         <= `TILE123.piton_pc_vld;
                  spc123_phy_pc_w          <= `TILE123.piton_pc;
                end
            end
    

            assign spc124_thread_id = 2'b00;
            assign spc124_rtl_pc = spc124_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(124*4)]   <= 1'b0;
                  active_thread[(124*4)+1] <= 1'b0;
                  active_thread[(124*4)+2] <= 1'b0;
                  active_thread[(124*4)+3] <= 1'b0;
                  spc124_inst_done         <= 0;
                  spc124_phy_pc_w          <= 0;
                end else begin
                  active_thread[(124*4)]   <= 1'b1;
                  active_thread[(124*4)+1] <= 1'b1;
                  active_thread[(124*4)+2] <= 1'b1;
                  active_thread[(124*4)+3] <= 1'b1;
                  spc124_inst_done         <= `TILE124.piton_pc_vld;
                  spc124_phy_pc_w          <= `TILE124.piton_pc;
                end
            end
    

            assign spc125_thread_id = 2'b00;
            assign spc125_rtl_pc = spc125_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(125*4)]   <= 1'b0;
                  active_thread[(125*4)+1] <= 1'b0;
                  active_thread[(125*4)+2] <= 1'b0;
                  active_thread[(125*4)+3] <= 1'b0;
                  spc125_inst_done         <= 0;
                  spc125_phy_pc_w          <= 0;
                end else begin
                  active_thread[(125*4)]   <= 1'b1;
                  active_thread[(125*4)+1] <= 1'b1;
                  active_thread[(125*4)+2] <= 1'b1;
                  active_thread[(125*4)+3] <= 1'b1;
                  spc125_inst_done         <= `TILE125.piton_pc_vld;
                  spc125_phy_pc_w          <= `TILE125.piton_pc;
                end
            end
    

            assign spc126_thread_id = 2'b00;
            assign spc126_rtl_pc = spc126_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(126*4)]   <= 1'b0;
                  active_thread[(126*4)+1] <= 1'b0;
                  active_thread[(126*4)+2] <= 1'b0;
                  active_thread[(126*4)+3] <= 1'b0;
                  spc126_inst_done         <= 0;
                  spc126_phy_pc_w          <= 0;
                end else begin
                  active_thread[(126*4)]   <= 1'b1;
                  active_thread[(126*4)+1] <= 1'b1;
                  active_thread[(126*4)+2] <= 1'b1;
                  active_thread[(126*4)+3] <= 1'b1;
                  spc126_inst_done         <= `TILE126.piton_pc_vld;
                  spc126_phy_pc_w          <= `TILE126.piton_pc;
                end
            end
    

            assign spc127_thread_id = 2'b00;
            assign spc127_rtl_pc = spc127_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(127*4)]   <= 1'b0;
                  active_thread[(127*4)+1] <= 1'b0;
                  active_thread[(127*4)+2] <= 1'b0;
                  active_thread[(127*4)+3] <= 1'b0;
                  spc127_inst_done         <= 0;
                  spc127_phy_pc_w          <= 0;
                end else begin
                  active_thread[(127*4)]   <= 1'b1;
                  active_thread[(127*4)+1] <= 1'b1;
                  active_thread[(127*4)+2] <= 1'b1;
                  active_thread[(127*4)+3] <= 1'b1;
                  spc127_inst_done         <= `TILE127.piton_pc_vld;
                  spc127_phy_pc_w          <= `TILE127.piton_pc;
                end
            end
    

            assign spc128_thread_id = 2'b00;
            assign spc128_rtl_pc = spc128_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(128*4)]   <= 1'b0;
                  active_thread[(128*4)+1] <= 1'b0;
                  active_thread[(128*4)+2] <= 1'b0;
                  active_thread[(128*4)+3] <= 1'b0;
                  spc128_inst_done         <= 0;
                  spc128_phy_pc_w          <= 0;
                end else begin
                  active_thread[(128*4)]   <= 1'b1;
                  active_thread[(128*4)+1] <= 1'b1;
                  active_thread[(128*4)+2] <= 1'b1;
                  active_thread[(128*4)+3] <= 1'b1;
                  spc128_inst_done         <= `TILE128.piton_pc_vld;
                  spc128_phy_pc_w          <= `TILE128.piton_pc;
                end
            end
    

            assign spc129_thread_id = 2'b00;
            assign spc129_rtl_pc = spc129_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(129*4)]   <= 1'b0;
                  active_thread[(129*4)+1] <= 1'b0;
                  active_thread[(129*4)+2] <= 1'b0;
                  active_thread[(129*4)+3] <= 1'b0;
                  spc129_inst_done         <= 0;
                  spc129_phy_pc_w          <= 0;
                end else begin
                  active_thread[(129*4)]   <= 1'b1;
                  active_thread[(129*4)+1] <= 1'b1;
                  active_thread[(129*4)+2] <= 1'b1;
                  active_thread[(129*4)+3] <= 1'b1;
                  spc129_inst_done         <= `TILE129.piton_pc_vld;
                  spc129_phy_pc_w          <= `TILE129.piton_pc;
                end
            end
    

            assign spc130_thread_id = 2'b00;
            assign spc130_rtl_pc = spc130_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(130*4)]   <= 1'b0;
                  active_thread[(130*4)+1] <= 1'b0;
                  active_thread[(130*4)+2] <= 1'b0;
                  active_thread[(130*4)+3] <= 1'b0;
                  spc130_inst_done         <= 0;
                  spc130_phy_pc_w          <= 0;
                end else begin
                  active_thread[(130*4)]   <= 1'b1;
                  active_thread[(130*4)+1] <= 1'b1;
                  active_thread[(130*4)+2] <= 1'b1;
                  active_thread[(130*4)+3] <= 1'b1;
                  spc130_inst_done         <= `TILE130.piton_pc_vld;
                  spc130_phy_pc_w          <= `TILE130.piton_pc;
                end
            end
    

            assign spc131_thread_id = 2'b00;
            assign spc131_rtl_pc = spc131_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(131*4)]   <= 1'b0;
                  active_thread[(131*4)+1] <= 1'b0;
                  active_thread[(131*4)+2] <= 1'b0;
                  active_thread[(131*4)+3] <= 1'b0;
                  spc131_inst_done         <= 0;
                  spc131_phy_pc_w          <= 0;
                end else begin
                  active_thread[(131*4)]   <= 1'b1;
                  active_thread[(131*4)+1] <= 1'b1;
                  active_thread[(131*4)+2] <= 1'b1;
                  active_thread[(131*4)+3] <= 1'b1;
                  spc131_inst_done         <= `TILE131.piton_pc_vld;
                  spc131_phy_pc_w          <= `TILE131.piton_pc;
                end
            end
    

            assign spc132_thread_id = 2'b00;
            assign spc132_rtl_pc = spc132_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(132*4)]   <= 1'b0;
                  active_thread[(132*4)+1] <= 1'b0;
                  active_thread[(132*4)+2] <= 1'b0;
                  active_thread[(132*4)+3] <= 1'b0;
                  spc132_inst_done         <= 0;
                  spc132_phy_pc_w          <= 0;
                end else begin
                  active_thread[(132*4)]   <= 1'b1;
                  active_thread[(132*4)+1] <= 1'b1;
                  active_thread[(132*4)+2] <= 1'b1;
                  active_thread[(132*4)+3] <= 1'b1;
                  spc132_inst_done         <= `TILE132.piton_pc_vld;
                  spc132_phy_pc_w          <= `TILE132.piton_pc;
                end
            end
    

            assign spc133_thread_id = 2'b00;
            assign spc133_rtl_pc = spc133_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(133*4)]   <= 1'b0;
                  active_thread[(133*4)+1] <= 1'b0;
                  active_thread[(133*4)+2] <= 1'b0;
                  active_thread[(133*4)+3] <= 1'b0;
                  spc133_inst_done         <= 0;
                  spc133_phy_pc_w          <= 0;
                end else begin
                  active_thread[(133*4)]   <= 1'b1;
                  active_thread[(133*4)+1] <= 1'b1;
                  active_thread[(133*4)+2] <= 1'b1;
                  active_thread[(133*4)+3] <= 1'b1;
                  spc133_inst_done         <= `TILE133.piton_pc_vld;
                  spc133_phy_pc_w          <= `TILE133.piton_pc;
                end
            end
    

            assign spc134_thread_id = 2'b00;
            assign spc134_rtl_pc = spc134_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(134*4)]   <= 1'b0;
                  active_thread[(134*4)+1] <= 1'b0;
                  active_thread[(134*4)+2] <= 1'b0;
                  active_thread[(134*4)+3] <= 1'b0;
                  spc134_inst_done         <= 0;
                  spc134_phy_pc_w          <= 0;
                end else begin
                  active_thread[(134*4)]   <= 1'b1;
                  active_thread[(134*4)+1] <= 1'b1;
                  active_thread[(134*4)+2] <= 1'b1;
                  active_thread[(134*4)+3] <= 1'b1;
                  spc134_inst_done         <= `TILE134.piton_pc_vld;
                  spc134_phy_pc_w          <= `TILE134.piton_pc;
                end
            end
    

            assign spc135_thread_id = 2'b00;
            assign spc135_rtl_pc = spc135_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(135*4)]   <= 1'b0;
                  active_thread[(135*4)+1] <= 1'b0;
                  active_thread[(135*4)+2] <= 1'b0;
                  active_thread[(135*4)+3] <= 1'b0;
                  spc135_inst_done         <= 0;
                  spc135_phy_pc_w          <= 0;
                end else begin
                  active_thread[(135*4)]   <= 1'b1;
                  active_thread[(135*4)+1] <= 1'b1;
                  active_thread[(135*4)+2] <= 1'b1;
                  active_thread[(135*4)+3] <= 1'b1;
                  spc135_inst_done         <= `TILE135.piton_pc_vld;
                  spc135_phy_pc_w          <= `TILE135.piton_pc;
                end
            end
    

            assign spc136_thread_id = 2'b00;
            assign spc136_rtl_pc = spc136_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(136*4)]   <= 1'b0;
                  active_thread[(136*4)+1] <= 1'b0;
                  active_thread[(136*4)+2] <= 1'b0;
                  active_thread[(136*4)+3] <= 1'b0;
                  spc136_inst_done         <= 0;
                  spc136_phy_pc_w          <= 0;
                end else begin
                  active_thread[(136*4)]   <= 1'b1;
                  active_thread[(136*4)+1] <= 1'b1;
                  active_thread[(136*4)+2] <= 1'b1;
                  active_thread[(136*4)+3] <= 1'b1;
                  spc136_inst_done         <= `TILE136.piton_pc_vld;
                  spc136_phy_pc_w          <= `TILE136.piton_pc;
                end
            end
    

            assign spc137_thread_id = 2'b00;
            assign spc137_rtl_pc = spc137_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(137*4)]   <= 1'b0;
                  active_thread[(137*4)+1] <= 1'b0;
                  active_thread[(137*4)+2] <= 1'b0;
                  active_thread[(137*4)+3] <= 1'b0;
                  spc137_inst_done         <= 0;
                  spc137_phy_pc_w          <= 0;
                end else begin
                  active_thread[(137*4)]   <= 1'b1;
                  active_thread[(137*4)+1] <= 1'b1;
                  active_thread[(137*4)+2] <= 1'b1;
                  active_thread[(137*4)+3] <= 1'b1;
                  spc137_inst_done         <= `TILE137.piton_pc_vld;
                  spc137_phy_pc_w          <= `TILE137.piton_pc;
                end
            end
    

            assign spc138_thread_id = 2'b00;
            assign spc138_rtl_pc = spc138_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(138*4)]   <= 1'b0;
                  active_thread[(138*4)+1] <= 1'b0;
                  active_thread[(138*4)+2] <= 1'b0;
                  active_thread[(138*4)+3] <= 1'b0;
                  spc138_inst_done         <= 0;
                  spc138_phy_pc_w          <= 0;
                end else begin
                  active_thread[(138*4)]   <= 1'b1;
                  active_thread[(138*4)+1] <= 1'b1;
                  active_thread[(138*4)+2] <= 1'b1;
                  active_thread[(138*4)+3] <= 1'b1;
                  spc138_inst_done         <= `TILE138.piton_pc_vld;
                  spc138_phy_pc_w          <= `TILE138.piton_pc;
                end
            end
    

            assign spc139_thread_id = 2'b00;
            assign spc139_rtl_pc = spc139_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(139*4)]   <= 1'b0;
                  active_thread[(139*4)+1] <= 1'b0;
                  active_thread[(139*4)+2] <= 1'b0;
                  active_thread[(139*4)+3] <= 1'b0;
                  spc139_inst_done         <= 0;
                  spc139_phy_pc_w          <= 0;
                end else begin
                  active_thread[(139*4)]   <= 1'b1;
                  active_thread[(139*4)+1] <= 1'b1;
                  active_thread[(139*4)+2] <= 1'b1;
                  active_thread[(139*4)+3] <= 1'b1;
                  spc139_inst_done         <= `TILE139.piton_pc_vld;
                  spc139_phy_pc_w          <= `TILE139.piton_pc;
                end
            end
    

            assign spc140_thread_id = 2'b00;
            assign spc140_rtl_pc = spc140_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(140*4)]   <= 1'b0;
                  active_thread[(140*4)+1] <= 1'b0;
                  active_thread[(140*4)+2] <= 1'b0;
                  active_thread[(140*4)+3] <= 1'b0;
                  spc140_inst_done         <= 0;
                  spc140_phy_pc_w          <= 0;
                end else begin
                  active_thread[(140*4)]   <= 1'b1;
                  active_thread[(140*4)+1] <= 1'b1;
                  active_thread[(140*4)+2] <= 1'b1;
                  active_thread[(140*4)+3] <= 1'b1;
                  spc140_inst_done         <= `TILE140.piton_pc_vld;
                  spc140_phy_pc_w          <= `TILE140.piton_pc;
                end
            end
    

            assign spc141_thread_id = 2'b00;
            assign spc141_rtl_pc = spc141_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(141*4)]   <= 1'b0;
                  active_thread[(141*4)+1] <= 1'b0;
                  active_thread[(141*4)+2] <= 1'b0;
                  active_thread[(141*4)+3] <= 1'b0;
                  spc141_inst_done         <= 0;
                  spc141_phy_pc_w          <= 0;
                end else begin
                  active_thread[(141*4)]   <= 1'b1;
                  active_thread[(141*4)+1] <= 1'b1;
                  active_thread[(141*4)+2] <= 1'b1;
                  active_thread[(141*4)+3] <= 1'b1;
                  spc141_inst_done         <= `TILE141.piton_pc_vld;
                  spc141_phy_pc_w          <= `TILE141.piton_pc;
                end
            end
    

            assign spc142_thread_id = 2'b00;
            assign spc142_rtl_pc = spc142_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(142*4)]   <= 1'b0;
                  active_thread[(142*4)+1] <= 1'b0;
                  active_thread[(142*4)+2] <= 1'b0;
                  active_thread[(142*4)+3] <= 1'b0;
                  spc142_inst_done         <= 0;
                  spc142_phy_pc_w          <= 0;
                end else begin
                  active_thread[(142*4)]   <= 1'b1;
                  active_thread[(142*4)+1] <= 1'b1;
                  active_thread[(142*4)+2] <= 1'b1;
                  active_thread[(142*4)+3] <= 1'b1;
                  spc142_inst_done         <= `TILE142.piton_pc_vld;
                  spc142_phy_pc_w          <= `TILE142.piton_pc;
                end
            end
    

            assign spc143_thread_id = 2'b00;
            assign spc143_rtl_pc = spc143_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(143*4)]   <= 1'b0;
                  active_thread[(143*4)+1] <= 1'b0;
                  active_thread[(143*4)+2] <= 1'b0;
                  active_thread[(143*4)+3] <= 1'b0;
                  spc143_inst_done         <= 0;
                  spc143_phy_pc_w          <= 0;
                end else begin
                  active_thread[(143*4)]   <= 1'b1;
                  active_thread[(143*4)+1] <= 1'b1;
                  active_thread[(143*4)+2] <= 1'b1;
                  active_thread[(143*4)+3] <= 1'b1;
                  spc143_inst_done         <= `TILE143.piton_pc_vld;
                  spc143_phy_pc_w          <= `TILE143.piton_pc;
                end
            end
    

            assign spc144_thread_id = 2'b00;
            assign spc144_rtl_pc = spc144_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(144*4)]   <= 1'b0;
                  active_thread[(144*4)+1] <= 1'b0;
                  active_thread[(144*4)+2] <= 1'b0;
                  active_thread[(144*4)+3] <= 1'b0;
                  spc144_inst_done         <= 0;
                  spc144_phy_pc_w          <= 0;
                end else begin
                  active_thread[(144*4)]   <= 1'b1;
                  active_thread[(144*4)+1] <= 1'b1;
                  active_thread[(144*4)+2] <= 1'b1;
                  active_thread[(144*4)+3] <= 1'b1;
                  spc144_inst_done         <= `TILE144.piton_pc_vld;
                  spc144_phy_pc_w          <= `TILE144.piton_pc;
                end
            end
    

            assign spc145_thread_id = 2'b00;
            assign spc145_rtl_pc = spc145_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(145*4)]   <= 1'b0;
                  active_thread[(145*4)+1] <= 1'b0;
                  active_thread[(145*4)+2] <= 1'b0;
                  active_thread[(145*4)+3] <= 1'b0;
                  spc145_inst_done         <= 0;
                  spc145_phy_pc_w          <= 0;
                end else begin
                  active_thread[(145*4)]   <= 1'b1;
                  active_thread[(145*4)+1] <= 1'b1;
                  active_thread[(145*4)+2] <= 1'b1;
                  active_thread[(145*4)+3] <= 1'b1;
                  spc145_inst_done         <= `TILE145.piton_pc_vld;
                  spc145_phy_pc_w          <= `TILE145.piton_pc;
                end
            end
    

            assign spc146_thread_id = 2'b00;
            assign spc146_rtl_pc = spc146_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(146*4)]   <= 1'b0;
                  active_thread[(146*4)+1] <= 1'b0;
                  active_thread[(146*4)+2] <= 1'b0;
                  active_thread[(146*4)+3] <= 1'b0;
                  spc146_inst_done         <= 0;
                  spc146_phy_pc_w          <= 0;
                end else begin
                  active_thread[(146*4)]   <= 1'b1;
                  active_thread[(146*4)+1] <= 1'b1;
                  active_thread[(146*4)+2] <= 1'b1;
                  active_thread[(146*4)+3] <= 1'b1;
                  spc146_inst_done         <= `TILE146.piton_pc_vld;
                  spc146_phy_pc_w          <= `TILE146.piton_pc;
                end
            end
    

            assign spc147_thread_id = 2'b00;
            assign spc147_rtl_pc = spc147_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(147*4)]   <= 1'b0;
                  active_thread[(147*4)+1] <= 1'b0;
                  active_thread[(147*4)+2] <= 1'b0;
                  active_thread[(147*4)+3] <= 1'b0;
                  spc147_inst_done         <= 0;
                  spc147_phy_pc_w          <= 0;
                end else begin
                  active_thread[(147*4)]   <= 1'b1;
                  active_thread[(147*4)+1] <= 1'b1;
                  active_thread[(147*4)+2] <= 1'b1;
                  active_thread[(147*4)+3] <= 1'b1;
                  spc147_inst_done         <= `TILE147.piton_pc_vld;
                  spc147_phy_pc_w          <= `TILE147.piton_pc;
                end
            end
    

            assign spc148_thread_id = 2'b00;
            assign spc148_rtl_pc = spc148_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(148*4)]   <= 1'b0;
                  active_thread[(148*4)+1] <= 1'b0;
                  active_thread[(148*4)+2] <= 1'b0;
                  active_thread[(148*4)+3] <= 1'b0;
                  spc148_inst_done         <= 0;
                  spc148_phy_pc_w          <= 0;
                end else begin
                  active_thread[(148*4)]   <= 1'b1;
                  active_thread[(148*4)+1] <= 1'b1;
                  active_thread[(148*4)+2] <= 1'b1;
                  active_thread[(148*4)+3] <= 1'b1;
                  spc148_inst_done         <= `TILE148.piton_pc_vld;
                  spc148_phy_pc_w          <= `TILE148.piton_pc;
                end
            end
    

            assign spc149_thread_id = 2'b00;
            assign spc149_rtl_pc = spc149_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(149*4)]   <= 1'b0;
                  active_thread[(149*4)+1] <= 1'b0;
                  active_thread[(149*4)+2] <= 1'b0;
                  active_thread[(149*4)+3] <= 1'b0;
                  spc149_inst_done         <= 0;
                  spc149_phy_pc_w          <= 0;
                end else begin
                  active_thread[(149*4)]   <= 1'b1;
                  active_thread[(149*4)+1] <= 1'b1;
                  active_thread[(149*4)+2] <= 1'b1;
                  active_thread[(149*4)+3] <= 1'b1;
                  spc149_inst_done         <= `TILE149.piton_pc_vld;
                  spc149_phy_pc_w          <= `TILE149.piton_pc;
                end
            end
    

            assign spc150_thread_id = 2'b00;
            assign spc150_rtl_pc = spc150_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(150*4)]   <= 1'b0;
                  active_thread[(150*4)+1] <= 1'b0;
                  active_thread[(150*4)+2] <= 1'b0;
                  active_thread[(150*4)+3] <= 1'b0;
                  spc150_inst_done         <= 0;
                  spc150_phy_pc_w          <= 0;
                end else begin
                  active_thread[(150*4)]   <= 1'b1;
                  active_thread[(150*4)+1] <= 1'b1;
                  active_thread[(150*4)+2] <= 1'b1;
                  active_thread[(150*4)+3] <= 1'b1;
                  spc150_inst_done         <= `TILE150.piton_pc_vld;
                  spc150_phy_pc_w          <= `TILE150.piton_pc;
                end
            end
    

            assign spc151_thread_id = 2'b00;
            assign spc151_rtl_pc = spc151_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(151*4)]   <= 1'b0;
                  active_thread[(151*4)+1] <= 1'b0;
                  active_thread[(151*4)+2] <= 1'b0;
                  active_thread[(151*4)+3] <= 1'b0;
                  spc151_inst_done         <= 0;
                  spc151_phy_pc_w          <= 0;
                end else begin
                  active_thread[(151*4)]   <= 1'b1;
                  active_thread[(151*4)+1] <= 1'b1;
                  active_thread[(151*4)+2] <= 1'b1;
                  active_thread[(151*4)+3] <= 1'b1;
                  spc151_inst_done         <= `TILE151.piton_pc_vld;
                  spc151_phy_pc_w          <= `TILE151.piton_pc;
                end
            end
    

            assign spc152_thread_id = 2'b00;
            assign spc152_rtl_pc = spc152_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(152*4)]   <= 1'b0;
                  active_thread[(152*4)+1] <= 1'b0;
                  active_thread[(152*4)+2] <= 1'b0;
                  active_thread[(152*4)+3] <= 1'b0;
                  spc152_inst_done         <= 0;
                  spc152_phy_pc_w          <= 0;
                end else begin
                  active_thread[(152*4)]   <= 1'b1;
                  active_thread[(152*4)+1] <= 1'b1;
                  active_thread[(152*4)+2] <= 1'b1;
                  active_thread[(152*4)+3] <= 1'b1;
                  spc152_inst_done         <= `TILE152.piton_pc_vld;
                  spc152_phy_pc_w          <= `TILE152.piton_pc;
                end
            end
    

            assign spc153_thread_id = 2'b00;
            assign spc153_rtl_pc = spc153_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(153*4)]   <= 1'b0;
                  active_thread[(153*4)+1] <= 1'b0;
                  active_thread[(153*4)+2] <= 1'b0;
                  active_thread[(153*4)+3] <= 1'b0;
                  spc153_inst_done         <= 0;
                  spc153_phy_pc_w          <= 0;
                end else begin
                  active_thread[(153*4)]   <= 1'b1;
                  active_thread[(153*4)+1] <= 1'b1;
                  active_thread[(153*4)+2] <= 1'b1;
                  active_thread[(153*4)+3] <= 1'b1;
                  spc153_inst_done         <= `TILE153.piton_pc_vld;
                  spc153_phy_pc_w          <= `TILE153.piton_pc;
                end
            end
    

            assign spc154_thread_id = 2'b00;
            assign spc154_rtl_pc = spc154_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(154*4)]   <= 1'b0;
                  active_thread[(154*4)+1] <= 1'b0;
                  active_thread[(154*4)+2] <= 1'b0;
                  active_thread[(154*4)+3] <= 1'b0;
                  spc154_inst_done         <= 0;
                  spc154_phy_pc_w          <= 0;
                end else begin
                  active_thread[(154*4)]   <= 1'b1;
                  active_thread[(154*4)+1] <= 1'b1;
                  active_thread[(154*4)+2] <= 1'b1;
                  active_thread[(154*4)+3] <= 1'b1;
                  spc154_inst_done         <= `TILE154.piton_pc_vld;
                  spc154_phy_pc_w          <= `TILE154.piton_pc;
                end
            end
    

            assign spc155_thread_id = 2'b00;
            assign spc155_rtl_pc = spc155_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(155*4)]   <= 1'b0;
                  active_thread[(155*4)+1] <= 1'b0;
                  active_thread[(155*4)+2] <= 1'b0;
                  active_thread[(155*4)+3] <= 1'b0;
                  spc155_inst_done         <= 0;
                  spc155_phy_pc_w          <= 0;
                end else begin
                  active_thread[(155*4)]   <= 1'b1;
                  active_thread[(155*4)+1] <= 1'b1;
                  active_thread[(155*4)+2] <= 1'b1;
                  active_thread[(155*4)+3] <= 1'b1;
                  spc155_inst_done         <= `TILE155.piton_pc_vld;
                  spc155_phy_pc_w          <= `TILE155.piton_pc;
                end
            end
    

            assign spc156_thread_id = 2'b00;
            assign spc156_rtl_pc = spc156_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(156*4)]   <= 1'b0;
                  active_thread[(156*4)+1] <= 1'b0;
                  active_thread[(156*4)+2] <= 1'b0;
                  active_thread[(156*4)+3] <= 1'b0;
                  spc156_inst_done         <= 0;
                  spc156_phy_pc_w          <= 0;
                end else begin
                  active_thread[(156*4)]   <= 1'b1;
                  active_thread[(156*4)+1] <= 1'b1;
                  active_thread[(156*4)+2] <= 1'b1;
                  active_thread[(156*4)+3] <= 1'b1;
                  spc156_inst_done         <= `TILE156.piton_pc_vld;
                  spc156_phy_pc_w          <= `TILE156.piton_pc;
                end
            end
    

            assign spc157_thread_id = 2'b00;
            assign spc157_rtl_pc = spc157_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(157*4)]   <= 1'b0;
                  active_thread[(157*4)+1] <= 1'b0;
                  active_thread[(157*4)+2] <= 1'b0;
                  active_thread[(157*4)+3] <= 1'b0;
                  spc157_inst_done         <= 0;
                  spc157_phy_pc_w          <= 0;
                end else begin
                  active_thread[(157*4)]   <= 1'b1;
                  active_thread[(157*4)+1] <= 1'b1;
                  active_thread[(157*4)+2] <= 1'b1;
                  active_thread[(157*4)+3] <= 1'b1;
                  spc157_inst_done         <= `TILE157.piton_pc_vld;
                  spc157_phy_pc_w          <= `TILE157.piton_pc;
                end
            end
    

            assign spc158_thread_id = 2'b00;
            assign spc158_rtl_pc = spc158_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(158*4)]   <= 1'b0;
                  active_thread[(158*4)+1] <= 1'b0;
                  active_thread[(158*4)+2] <= 1'b0;
                  active_thread[(158*4)+3] <= 1'b0;
                  spc158_inst_done         <= 0;
                  spc158_phy_pc_w          <= 0;
                end else begin
                  active_thread[(158*4)]   <= 1'b1;
                  active_thread[(158*4)+1] <= 1'b1;
                  active_thread[(158*4)+2] <= 1'b1;
                  active_thread[(158*4)+3] <= 1'b1;
                  spc158_inst_done         <= `TILE158.piton_pc_vld;
                  spc158_phy_pc_w          <= `TILE158.piton_pc;
                end
            end
    

            assign spc159_thread_id = 2'b00;
            assign spc159_rtl_pc = spc159_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(159*4)]   <= 1'b0;
                  active_thread[(159*4)+1] <= 1'b0;
                  active_thread[(159*4)+2] <= 1'b0;
                  active_thread[(159*4)+3] <= 1'b0;
                  spc159_inst_done         <= 0;
                  spc159_phy_pc_w          <= 0;
                end else begin
                  active_thread[(159*4)]   <= 1'b1;
                  active_thread[(159*4)+1] <= 1'b1;
                  active_thread[(159*4)+2] <= 1'b1;
                  active_thread[(159*4)+3] <= 1'b1;
                  spc159_inst_done         <= `TILE159.piton_pc_vld;
                  spc159_phy_pc_w          <= `TILE159.piton_pc;
                end
            end
    

            assign spc160_thread_id = 2'b00;
            assign spc160_rtl_pc = spc160_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(160*4)]   <= 1'b0;
                  active_thread[(160*4)+1] <= 1'b0;
                  active_thread[(160*4)+2] <= 1'b0;
                  active_thread[(160*4)+3] <= 1'b0;
                  spc160_inst_done         <= 0;
                  spc160_phy_pc_w          <= 0;
                end else begin
                  active_thread[(160*4)]   <= 1'b1;
                  active_thread[(160*4)+1] <= 1'b1;
                  active_thread[(160*4)+2] <= 1'b1;
                  active_thread[(160*4)+3] <= 1'b1;
                  spc160_inst_done         <= `TILE160.piton_pc_vld;
                  spc160_phy_pc_w          <= `TILE160.piton_pc;
                end
            end
    

            assign spc161_thread_id = 2'b00;
            assign spc161_rtl_pc = spc161_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(161*4)]   <= 1'b0;
                  active_thread[(161*4)+1] <= 1'b0;
                  active_thread[(161*4)+2] <= 1'b0;
                  active_thread[(161*4)+3] <= 1'b0;
                  spc161_inst_done         <= 0;
                  spc161_phy_pc_w          <= 0;
                end else begin
                  active_thread[(161*4)]   <= 1'b1;
                  active_thread[(161*4)+1] <= 1'b1;
                  active_thread[(161*4)+2] <= 1'b1;
                  active_thread[(161*4)+3] <= 1'b1;
                  spc161_inst_done         <= `TILE161.piton_pc_vld;
                  spc161_phy_pc_w          <= `TILE161.piton_pc;
                end
            end
    

            assign spc162_thread_id = 2'b00;
            assign spc162_rtl_pc = spc162_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(162*4)]   <= 1'b0;
                  active_thread[(162*4)+1] <= 1'b0;
                  active_thread[(162*4)+2] <= 1'b0;
                  active_thread[(162*4)+3] <= 1'b0;
                  spc162_inst_done         <= 0;
                  spc162_phy_pc_w          <= 0;
                end else begin
                  active_thread[(162*4)]   <= 1'b1;
                  active_thread[(162*4)+1] <= 1'b1;
                  active_thread[(162*4)+2] <= 1'b1;
                  active_thread[(162*4)+3] <= 1'b1;
                  spc162_inst_done         <= `TILE162.piton_pc_vld;
                  spc162_phy_pc_w          <= `TILE162.piton_pc;
                end
            end
    

            assign spc163_thread_id = 2'b00;
            assign spc163_rtl_pc = spc163_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(163*4)]   <= 1'b0;
                  active_thread[(163*4)+1] <= 1'b0;
                  active_thread[(163*4)+2] <= 1'b0;
                  active_thread[(163*4)+3] <= 1'b0;
                  spc163_inst_done         <= 0;
                  spc163_phy_pc_w          <= 0;
                end else begin
                  active_thread[(163*4)]   <= 1'b1;
                  active_thread[(163*4)+1] <= 1'b1;
                  active_thread[(163*4)+2] <= 1'b1;
                  active_thread[(163*4)+3] <= 1'b1;
                  spc163_inst_done         <= `TILE163.piton_pc_vld;
                  spc163_phy_pc_w          <= `TILE163.piton_pc;
                end
            end
    

            assign spc164_thread_id = 2'b00;
            assign spc164_rtl_pc = spc164_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(164*4)]   <= 1'b0;
                  active_thread[(164*4)+1] <= 1'b0;
                  active_thread[(164*4)+2] <= 1'b0;
                  active_thread[(164*4)+3] <= 1'b0;
                  spc164_inst_done         <= 0;
                  spc164_phy_pc_w          <= 0;
                end else begin
                  active_thread[(164*4)]   <= 1'b1;
                  active_thread[(164*4)+1] <= 1'b1;
                  active_thread[(164*4)+2] <= 1'b1;
                  active_thread[(164*4)+3] <= 1'b1;
                  spc164_inst_done         <= `TILE164.piton_pc_vld;
                  spc164_phy_pc_w          <= `TILE164.piton_pc;
                end
            end
    

            assign spc165_thread_id = 2'b00;
            assign spc165_rtl_pc = spc165_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(165*4)]   <= 1'b0;
                  active_thread[(165*4)+1] <= 1'b0;
                  active_thread[(165*4)+2] <= 1'b0;
                  active_thread[(165*4)+3] <= 1'b0;
                  spc165_inst_done         <= 0;
                  spc165_phy_pc_w          <= 0;
                end else begin
                  active_thread[(165*4)]   <= 1'b1;
                  active_thread[(165*4)+1] <= 1'b1;
                  active_thread[(165*4)+2] <= 1'b1;
                  active_thread[(165*4)+3] <= 1'b1;
                  spc165_inst_done         <= `TILE165.piton_pc_vld;
                  spc165_phy_pc_w          <= `TILE165.piton_pc;
                end
            end
    

            assign spc166_thread_id = 2'b00;
            assign spc166_rtl_pc = spc166_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(166*4)]   <= 1'b0;
                  active_thread[(166*4)+1] <= 1'b0;
                  active_thread[(166*4)+2] <= 1'b0;
                  active_thread[(166*4)+3] <= 1'b0;
                  spc166_inst_done         <= 0;
                  spc166_phy_pc_w          <= 0;
                end else begin
                  active_thread[(166*4)]   <= 1'b1;
                  active_thread[(166*4)+1] <= 1'b1;
                  active_thread[(166*4)+2] <= 1'b1;
                  active_thread[(166*4)+3] <= 1'b1;
                  spc166_inst_done         <= `TILE166.piton_pc_vld;
                  spc166_phy_pc_w          <= `TILE166.piton_pc;
                end
            end
    

            assign spc167_thread_id = 2'b00;
            assign spc167_rtl_pc = spc167_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(167*4)]   <= 1'b0;
                  active_thread[(167*4)+1] <= 1'b0;
                  active_thread[(167*4)+2] <= 1'b0;
                  active_thread[(167*4)+3] <= 1'b0;
                  spc167_inst_done         <= 0;
                  spc167_phy_pc_w          <= 0;
                end else begin
                  active_thread[(167*4)]   <= 1'b1;
                  active_thread[(167*4)+1] <= 1'b1;
                  active_thread[(167*4)+2] <= 1'b1;
                  active_thread[(167*4)+3] <= 1'b1;
                  spc167_inst_done         <= `TILE167.piton_pc_vld;
                  spc167_phy_pc_w          <= `TILE167.piton_pc;
                end
            end
    

            assign spc168_thread_id = 2'b00;
            assign spc168_rtl_pc = spc168_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(168*4)]   <= 1'b0;
                  active_thread[(168*4)+1] <= 1'b0;
                  active_thread[(168*4)+2] <= 1'b0;
                  active_thread[(168*4)+3] <= 1'b0;
                  spc168_inst_done         <= 0;
                  spc168_phy_pc_w          <= 0;
                end else begin
                  active_thread[(168*4)]   <= 1'b1;
                  active_thread[(168*4)+1] <= 1'b1;
                  active_thread[(168*4)+2] <= 1'b1;
                  active_thread[(168*4)+3] <= 1'b1;
                  spc168_inst_done         <= `TILE168.piton_pc_vld;
                  spc168_phy_pc_w          <= `TILE168.piton_pc;
                end
            end
    

            assign spc169_thread_id = 2'b00;
            assign spc169_rtl_pc = spc169_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(169*4)]   <= 1'b0;
                  active_thread[(169*4)+1] <= 1'b0;
                  active_thread[(169*4)+2] <= 1'b0;
                  active_thread[(169*4)+3] <= 1'b0;
                  spc169_inst_done         <= 0;
                  spc169_phy_pc_w          <= 0;
                end else begin
                  active_thread[(169*4)]   <= 1'b1;
                  active_thread[(169*4)+1] <= 1'b1;
                  active_thread[(169*4)+2] <= 1'b1;
                  active_thread[(169*4)+3] <= 1'b1;
                  spc169_inst_done         <= `TILE169.piton_pc_vld;
                  spc169_phy_pc_w          <= `TILE169.piton_pc;
                end
            end
    

            assign spc170_thread_id = 2'b00;
            assign spc170_rtl_pc = spc170_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(170*4)]   <= 1'b0;
                  active_thread[(170*4)+1] <= 1'b0;
                  active_thread[(170*4)+2] <= 1'b0;
                  active_thread[(170*4)+3] <= 1'b0;
                  spc170_inst_done         <= 0;
                  spc170_phy_pc_w          <= 0;
                end else begin
                  active_thread[(170*4)]   <= 1'b1;
                  active_thread[(170*4)+1] <= 1'b1;
                  active_thread[(170*4)+2] <= 1'b1;
                  active_thread[(170*4)+3] <= 1'b1;
                  spc170_inst_done         <= `TILE170.piton_pc_vld;
                  spc170_phy_pc_w          <= `TILE170.piton_pc;
                end
            end
    

            assign spc171_thread_id = 2'b00;
            assign spc171_rtl_pc = spc171_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(171*4)]   <= 1'b0;
                  active_thread[(171*4)+1] <= 1'b0;
                  active_thread[(171*4)+2] <= 1'b0;
                  active_thread[(171*4)+3] <= 1'b0;
                  spc171_inst_done         <= 0;
                  spc171_phy_pc_w          <= 0;
                end else begin
                  active_thread[(171*4)]   <= 1'b1;
                  active_thread[(171*4)+1] <= 1'b1;
                  active_thread[(171*4)+2] <= 1'b1;
                  active_thread[(171*4)+3] <= 1'b1;
                  spc171_inst_done         <= `TILE171.piton_pc_vld;
                  spc171_phy_pc_w          <= `TILE171.piton_pc;
                end
            end
    

            assign spc172_thread_id = 2'b00;
            assign spc172_rtl_pc = spc172_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(172*4)]   <= 1'b0;
                  active_thread[(172*4)+1] <= 1'b0;
                  active_thread[(172*4)+2] <= 1'b0;
                  active_thread[(172*4)+3] <= 1'b0;
                  spc172_inst_done         <= 0;
                  spc172_phy_pc_w          <= 0;
                end else begin
                  active_thread[(172*4)]   <= 1'b1;
                  active_thread[(172*4)+1] <= 1'b1;
                  active_thread[(172*4)+2] <= 1'b1;
                  active_thread[(172*4)+3] <= 1'b1;
                  spc172_inst_done         <= `TILE172.piton_pc_vld;
                  spc172_phy_pc_w          <= `TILE172.piton_pc;
                end
            end
    

            assign spc173_thread_id = 2'b00;
            assign spc173_rtl_pc = spc173_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(173*4)]   <= 1'b0;
                  active_thread[(173*4)+1] <= 1'b0;
                  active_thread[(173*4)+2] <= 1'b0;
                  active_thread[(173*4)+3] <= 1'b0;
                  spc173_inst_done         <= 0;
                  spc173_phy_pc_w          <= 0;
                end else begin
                  active_thread[(173*4)]   <= 1'b1;
                  active_thread[(173*4)+1] <= 1'b1;
                  active_thread[(173*4)+2] <= 1'b1;
                  active_thread[(173*4)+3] <= 1'b1;
                  spc173_inst_done         <= `TILE173.piton_pc_vld;
                  spc173_phy_pc_w          <= `TILE173.piton_pc;
                end
            end
    

            assign spc174_thread_id = 2'b00;
            assign spc174_rtl_pc = spc174_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(174*4)]   <= 1'b0;
                  active_thread[(174*4)+1] <= 1'b0;
                  active_thread[(174*4)+2] <= 1'b0;
                  active_thread[(174*4)+3] <= 1'b0;
                  spc174_inst_done         <= 0;
                  spc174_phy_pc_w          <= 0;
                end else begin
                  active_thread[(174*4)]   <= 1'b1;
                  active_thread[(174*4)+1] <= 1'b1;
                  active_thread[(174*4)+2] <= 1'b1;
                  active_thread[(174*4)+3] <= 1'b1;
                  spc174_inst_done         <= `TILE174.piton_pc_vld;
                  spc174_phy_pc_w          <= `TILE174.piton_pc;
                end
            end
    

            assign spc175_thread_id = 2'b00;
            assign spc175_rtl_pc = spc175_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(175*4)]   <= 1'b0;
                  active_thread[(175*4)+1] <= 1'b0;
                  active_thread[(175*4)+2] <= 1'b0;
                  active_thread[(175*4)+3] <= 1'b0;
                  spc175_inst_done         <= 0;
                  spc175_phy_pc_w          <= 0;
                end else begin
                  active_thread[(175*4)]   <= 1'b1;
                  active_thread[(175*4)+1] <= 1'b1;
                  active_thread[(175*4)+2] <= 1'b1;
                  active_thread[(175*4)+3] <= 1'b1;
                  spc175_inst_done         <= `TILE175.piton_pc_vld;
                  spc175_phy_pc_w          <= `TILE175.piton_pc;
                end
            end
    

            assign spc176_thread_id = 2'b00;
            assign spc176_rtl_pc = spc176_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(176*4)]   <= 1'b0;
                  active_thread[(176*4)+1] <= 1'b0;
                  active_thread[(176*4)+2] <= 1'b0;
                  active_thread[(176*4)+3] <= 1'b0;
                  spc176_inst_done         <= 0;
                  spc176_phy_pc_w          <= 0;
                end else begin
                  active_thread[(176*4)]   <= 1'b1;
                  active_thread[(176*4)+1] <= 1'b1;
                  active_thread[(176*4)+2] <= 1'b1;
                  active_thread[(176*4)+3] <= 1'b1;
                  spc176_inst_done         <= `TILE176.piton_pc_vld;
                  spc176_phy_pc_w          <= `TILE176.piton_pc;
                end
            end
    

            assign spc177_thread_id = 2'b00;
            assign spc177_rtl_pc = spc177_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(177*4)]   <= 1'b0;
                  active_thread[(177*4)+1] <= 1'b0;
                  active_thread[(177*4)+2] <= 1'b0;
                  active_thread[(177*4)+3] <= 1'b0;
                  spc177_inst_done         <= 0;
                  spc177_phy_pc_w          <= 0;
                end else begin
                  active_thread[(177*4)]   <= 1'b1;
                  active_thread[(177*4)+1] <= 1'b1;
                  active_thread[(177*4)+2] <= 1'b1;
                  active_thread[(177*4)+3] <= 1'b1;
                  spc177_inst_done         <= `TILE177.piton_pc_vld;
                  spc177_phy_pc_w          <= `TILE177.piton_pc;
                end
            end
    

            assign spc178_thread_id = 2'b00;
            assign spc178_rtl_pc = spc178_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(178*4)]   <= 1'b0;
                  active_thread[(178*4)+1] <= 1'b0;
                  active_thread[(178*4)+2] <= 1'b0;
                  active_thread[(178*4)+3] <= 1'b0;
                  spc178_inst_done         <= 0;
                  spc178_phy_pc_w          <= 0;
                end else begin
                  active_thread[(178*4)]   <= 1'b1;
                  active_thread[(178*4)+1] <= 1'b1;
                  active_thread[(178*4)+2] <= 1'b1;
                  active_thread[(178*4)+3] <= 1'b1;
                  spc178_inst_done         <= `TILE178.piton_pc_vld;
                  spc178_phy_pc_w          <= `TILE178.piton_pc;
                end
            end
    

            assign spc179_thread_id = 2'b00;
            assign spc179_rtl_pc = spc179_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(179*4)]   <= 1'b0;
                  active_thread[(179*4)+1] <= 1'b0;
                  active_thread[(179*4)+2] <= 1'b0;
                  active_thread[(179*4)+3] <= 1'b0;
                  spc179_inst_done         <= 0;
                  spc179_phy_pc_w          <= 0;
                end else begin
                  active_thread[(179*4)]   <= 1'b1;
                  active_thread[(179*4)+1] <= 1'b1;
                  active_thread[(179*4)+2] <= 1'b1;
                  active_thread[(179*4)+3] <= 1'b1;
                  spc179_inst_done         <= `TILE179.piton_pc_vld;
                  spc179_phy_pc_w          <= `TILE179.piton_pc;
                end
            end
    

            assign spc180_thread_id = 2'b00;
            assign spc180_rtl_pc = spc180_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(180*4)]   <= 1'b0;
                  active_thread[(180*4)+1] <= 1'b0;
                  active_thread[(180*4)+2] <= 1'b0;
                  active_thread[(180*4)+3] <= 1'b0;
                  spc180_inst_done         <= 0;
                  spc180_phy_pc_w          <= 0;
                end else begin
                  active_thread[(180*4)]   <= 1'b1;
                  active_thread[(180*4)+1] <= 1'b1;
                  active_thread[(180*4)+2] <= 1'b1;
                  active_thread[(180*4)+3] <= 1'b1;
                  spc180_inst_done         <= `TILE180.piton_pc_vld;
                  spc180_phy_pc_w          <= `TILE180.piton_pc;
                end
            end
    

            assign spc181_thread_id = 2'b00;
            assign spc181_rtl_pc = spc181_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(181*4)]   <= 1'b0;
                  active_thread[(181*4)+1] <= 1'b0;
                  active_thread[(181*4)+2] <= 1'b0;
                  active_thread[(181*4)+3] <= 1'b0;
                  spc181_inst_done         <= 0;
                  spc181_phy_pc_w          <= 0;
                end else begin
                  active_thread[(181*4)]   <= 1'b1;
                  active_thread[(181*4)+1] <= 1'b1;
                  active_thread[(181*4)+2] <= 1'b1;
                  active_thread[(181*4)+3] <= 1'b1;
                  spc181_inst_done         <= `TILE181.piton_pc_vld;
                  spc181_phy_pc_w          <= `TILE181.piton_pc;
                end
            end
    

            assign spc182_thread_id = 2'b00;
            assign spc182_rtl_pc = spc182_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(182*4)]   <= 1'b0;
                  active_thread[(182*4)+1] <= 1'b0;
                  active_thread[(182*4)+2] <= 1'b0;
                  active_thread[(182*4)+3] <= 1'b0;
                  spc182_inst_done         <= 0;
                  spc182_phy_pc_w          <= 0;
                end else begin
                  active_thread[(182*4)]   <= 1'b1;
                  active_thread[(182*4)+1] <= 1'b1;
                  active_thread[(182*4)+2] <= 1'b1;
                  active_thread[(182*4)+3] <= 1'b1;
                  spc182_inst_done         <= `TILE182.piton_pc_vld;
                  spc182_phy_pc_w          <= `TILE182.piton_pc;
                end
            end
    

            assign spc183_thread_id = 2'b00;
            assign spc183_rtl_pc = spc183_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(183*4)]   <= 1'b0;
                  active_thread[(183*4)+1] <= 1'b0;
                  active_thread[(183*4)+2] <= 1'b0;
                  active_thread[(183*4)+3] <= 1'b0;
                  spc183_inst_done         <= 0;
                  spc183_phy_pc_w          <= 0;
                end else begin
                  active_thread[(183*4)]   <= 1'b1;
                  active_thread[(183*4)+1] <= 1'b1;
                  active_thread[(183*4)+2] <= 1'b1;
                  active_thread[(183*4)+3] <= 1'b1;
                  spc183_inst_done         <= `TILE183.piton_pc_vld;
                  spc183_phy_pc_w          <= `TILE183.piton_pc;
                end
            end
    

            assign spc184_thread_id = 2'b00;
            assign spc184_rtl_pc = spc184_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(184*4)]   <= 1'b0;
                  active_thread[(184*4)+1] <= 1'b0;
                  active_thread[(184*4)+2] <= 1'b0;
                  active_thread[(184*4)+3] <= 1'b0;
                  spc184_inst_done         <= 0;
                  spc184_phy_pc_w          <= 0;
                end else begin
                  active_thread[(184*4)]   <= 1'b1;
                  active_thread[(184*4)+1] <= 1'b1;
                  active_thread[(184*4)+2] <= 1'b1;
                  active_thread[(184*4)+3] <= 1'b1;
                  spc184_inst_done         <= `TILE184.piton_pc_vld;
                  spc184_phy_pc_w          <= `TILE184.piton_pc;
                end
            end
    

            assign spc185_thread_id = 2'b00;
            assign spc185_rtl_pc = spc185_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(185*4)]   <= 1'b0;
                  active_thread[(185*4)+1] <= 1'b0;
                  active_thread[(185*4)+2] <= 1'b0;
                  active_thread[(185*4)+3] <= 1'b0;
                  spc185_inst_done         <= 0;
                  spc185_phy_pc_w          <= 0;
                end else begin
                  active_thread[(185*4)]   <= 1'b1;
                  active_thread[(185*4)+1] <= 1'b1;
                  active_thread[(185*4)+2] <= 1'b1;
                  active_thread[(185*4)+3] <= 1'b1;
                  spc185_inst_done         <= `TILE185.piton_pc_vld;
                  spc185_phy_pc_w          <= `TILE185.piton_pc;
                end
            end
    

            assign spc186_thread_id = 2'b00;
            assign spc186_rtl_pc = spc186_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(186*4)]   <= 1'b0;
                  active_thread[(186*4)+1] <= 1'b0;
                  active_thread[(186*4)+2] <= 1'b0;
                  active_thread[(186*4)+3] <= 1'b0;
                  spc186_inst_done         <= 0;
                  spc186_phy_pc_w          <= 0;
                end else begin
                  active_thread[(186*4)]   <= 1'b1;
                  active_thread[(186*4)+1] <= 1'b1;
                  active_thread[(186*4)+2] <= 1'b1;
                  active_thread[(186*4)+3] <= 1'b1;
                  spc186_inst_done         <= `TILE186.piton_pc_vld;
                  spc186_phy_pc_w          <= `TILE186.piton_pc;
                end
            end
    

            assign spc187_thread_id = 2'b00;
            assign spc187_rtl_pc = spc187_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(187*4)]   <= 1'b0;
                  active_thread[(187*4)+1] <= 1'b0;
                  active_thread[(187*4)+2] <= 1'b0;
                  active_thread[(187*4)+3] <= 1'b0;
                  spc187_inst_done         <= 0;
                  spc187_phy_pc_w          <= 0;
                end else begin
                  active_thread[(187*4)]   <= 1'b1;
                  active_thread[(187*4)+1] <= 1'b1;
                  active_thread[(187*4)+2] <= 1'b1;
                  active_thread[(187*4)+3] <= 1'b1;
                  spc187_inst_done         <= `TILE187.piton_pc_vld;
                  spc187_phy_pc_w          <= `TILE187.piton_pc;
                end
            end
    

            assign spc188_thread_id = 2'b00;
            assign spc188_rtl_pc = spc188_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(188*4)]   <= 1'b0;
                  active_thread[(188*4)+1] <= 1'b0;
                  active_thread[(188*4)+2] <= 1'b0;
                  active_thread[(188*4)+3] <= 1'b0;
                  spc188_inst_done         <= 0;
                  spc188_phy_pc_w          <= 0;
                end else begin
                  active_thread[(188*4)]   <= 1'b1;
                  active_thread[(188*4)+1] <= 1'b1;
                  active_thread[(188*4)+2] <= 1'b1;
                  active_thread[(188*4)+3] <= 1'b1;
                  spc188_inst_done         <= `TILE188.piton_pc_vld;
                  spc188_phy_pc_w          <= `TILE188.piton_pc;
                end
            end
    

            assign spc189_thread_id = 2'b00;
            assign spc189_rtl_pc = spc189_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(189*4)]   <= 1'b0;
                  active_thread[(189*4)+1] <= 1'b0;
                  active_thread[(189*4)+2] <= 1'b0;
                  active_thread[(189*4)+3] <= 1'b0;
                  spc189_inst_done         <= 0;
                  spc189_phy_pc_w          <= 0;
                end else begin
                  active_thread[(189*4)]   <= 1'b1;
                  active_thread[(189*4)+1] <= 1'b1;
                  active_thread[(189*4)+2] <= 1'b1;
                  active_thread[(189*4)+3] <= 1'b1;
                  spc189_inst_done         <= `TILE189.piton_pc_vld;
                  spc189_phy_pc_w          <= `TILE189.piton_pc;
                end
            end
    

            assign spc190_thread_id = 2'b00;
            assign spc190_rtl_pc = spc190_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(190*4)]   <= 1'b0;
                  active_thread[(190*4)+1] <= 1'b0;
                  active_thread[(190*4)+2] <= 1'b0;
                  active_thread[(190*4)+3] <= 1'b0;
                  spc190_inst_done         <= 0;
                  spc190_phy_pc_w          <= 0;
                end else begin
                  active_thread[(190*4)]   <= 1'b1;
                  active_thread[(190*4)+1] <= 1'b1;
                  active_thread[(190*4)+2] <= 1'b1;
                  active_thread[(190*4)+3] <= 1'b1;
                  spc190_inst_done         <= `TILE190.piton_pc_vld;
                  spc190_phy_pc_w          <= `TILE190.piton_pc;
                end
            end
    

            assign spc191_thread_id = 2'b00;
            assign spc191_rtl_pc = spc191_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(191*4)]   <= 1'b0;
                  active_thread[(191*4)+1] <= 1'b0;
                  active_thread[(191*4)+2] <= 1'b0;
                  active_thread[(191*4)+3] <= 1'b0;
                  spc191_inst_done         <= 0;
                  spc191_phy_pc_w          <= 0;
                end else begin
                  active_thread[(191*4)]   <= 1'b1;
                  active_thread[(191*4)+1] <= 1'b1;
                  active_thread[(191*4)+2] <= 1'b1;
                  active_thread[(191*4)+3] <= 1'b1;
                  spc191_inst_done         <= `TILE191.piton_pc_vld;
                  spc191_phy_pc_w          <= `TILE191.piton_pc;
                end
            end
    

            assign spc192_thread_id = 2'b00;
            assign spc192_rtl_pc = spc192_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(192*4)]   <= 1'b0;
                  active_thread[(192*4)+1] <= 1'b0;
                  active_thread[(192*4)+2] <= 1'b0;
                  active_thread[(192*4)+3] <= 1'b0;
                  spc192_inst_done         <= 0;
                  spc192_phy_pc_w          <= 0;
                end else begin
                  active_thread[(192*4)]   <= 1'b1;
                  active_thread[(192*4)+1] <= 1'b1;
                  active_thread[(192*4)+2] <= 1'b1;
                  active_thread[(192*4)+3] <= 1'b1;
                  spc192_inst_done         <= `TILE192.piton_pc_vld;
                  spc192_phy_pc_w          <= `TILE192.piton_pc;
                end
            end
    

            assign spc193_thread_id = 2'b00;
            assign spc193_rtl_pc = spc193_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(193*4)]   <= 1'b0;
                  active_thread[(193*4)+1] <= 1'b0;
                  active_thread[(193*4)+2] <= 1'b0;
                  active_thread[(193*4)+3] <= 1'b0;
                  spc193_inst_done         <= 0;
                  spc193_phy_pc_w          <= 0;
                end else begin
                  active_thread[(193*4)]   <= 1'b1;
                  active_thread[(193*4)+1] <= 1'b1;
                  active_thread[(193*4)+2] <= 1'b1;
                  active_thread[(193*4)+3] <= 1'b1;
                  spc193_inst_done         <= `TILE193.piton_pc_vld;
                  spc193_phy_pc_w          <= `TILE193.piton_pc;
                end
            end
    

            assign spc194_thread_id = 2'b00;
            assign spc194_rtl_pc = spc194_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(194*4)]   <= 1'b0;
                  active_thread[(194*4)+1] <= 1'b0;
                  active_thread[(194*4)+2] <= 1'b0;
                  active_thread[(194*4)+3] <= 1'b0;
                  spc194_inst_done         <= 0;
                  spc194_phy_pc_w          <= 0;
                end else begin
                  active_thread[(194*4)]   <= 1'b1;
                  active_thread[(194*4)+1] <= 1'b1;
                  active_thread[(194*4)+2] <= 1'b1;
                  active_thread[(194*4)+3] <= 1'b1;
                  spc194_inst_done         <= `TILE194.piton_pc_vld;
                  spc194_phy_pc_w          <= `TILE194.piton_pc;
                end
            end
    

            assign spc195_thread_id = 2'b00;
            assign spc195_rtl_pc = spc195_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(195*4)]   <= 1'b0;
                  active_thread[(195*4)+1] <= 1'b0;
                  active_thread[(195*4)+2] <= 1'b0;
                  active_thread[(195*4)+3] <= 1'b0;
                  spc195_inst_done         <= 0;
                  spc195_phy_pc_w          <= 0;
                end else begin
                  active_thread[(195*4)]   <= 1'b1;
                  active_thread[(195*4)+1] <= 1'b1;
                  active_thread[(195*4)+2] <= 1'b1;
                  active_thread[(195*4)+3] <= 1'b1;
                  spc195_inst_done         <= `TILE195.piton_pc_vld;
                  spc195_phy_pc_w          <= `TILE195.piton_pc;
                end
            end
    

            assign spc196_thread_id = 2'b00;
            assign spc196_rtl_pc = spc196_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(196*4)]   <= 1'b0;
                  active_thread[(196*4)+1] <= 1'b0;
                  active_thread[(196*4)+2] <= 1'b0;
                  active_thread[(196*4)+3] <= 1'b0;
                  spc196_inst_done         <= 0;
                  spc196_phy_pc_w          <= 0;
                end else begin
                  active_thread[(196*4)]   <= 1'b1;
                  active_thread[(196*4)+1] <= 1'b1;
                  active_thread[(196*4)+2] <= 1'b1;
                  active_thread[(196*4)+3] <= 1'b1;
                  spc196_inst_done         <= `TILE196.piton_pc_vld;
                  spc196_phy_pc_w          <= `TILE196.piton_pc;
                end
            end
    

            assign spc197_thread_id = 2'b00;
            assign spc197_rtl_pc = spc197_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(197*4)]   <= 1'b0;
                  active_thread[(197*4)+1] <= 1'b0;
                  active_thread[(197*4)+2] <= 1'b0;
                  active_thread[(197*4)+3] <= 1'b0;
                  spc197_inst_done         <= 0;
                  spc197_phy_pc_w          <= 0;
                end else begin
                  active_thread[(197*4)]   <= 1'b1;
                  active_thread[(197*4)+1] <= 1'b1;
                  active_thread[(197*4)+2] <= 1'b1;
                  active_thread[(197*4)+3] <= 1'b1;
                  spc197_inst_done         <= `TILE197.piton_pc_vld;
                  spc197_phy_pc_w          <= `TILE197.piton_pc;
                end
            end
    

            assign spc198_thread_id = 2'b00;
            assign spc198_rtl_pc = spc198_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(198*4)]   <= 1'b0;
                  active_thread[(198*4)+1] <= 1'b0;
                  active_thread[(198*4)+2] <= 1'b0;
                  active_thread[(198*4)+3] <= 1'b0;
                  spc198_inst_done         <= 0;
                  spc198_phy_pc_w          <= 0;
                end else begin
                  active_thread[(198*4)]   <= 1'b1;
                  active_thread[(198*4)+1] <= 1'b1;
                  active_thread[(198*4)+2] <= 1'b1;
                  active_thread[(198*4)+3] <= 1'b1;
                  spc198_inst_done         <= `TILE198.piton_pc_vld;
                  spc198_phy_pc_w          <= `TILE198.piton_pc;
                end
            end
    

            assign spc199_thread_id = 2'b00;
            assign spc199_rtl_pc = spc199_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(199*4)]   <= 1'b0;
                  active_thread[(199*4)+1] <= 1'b0;
                  active_thread[(199*4)+2] <= 1'b0;
                  active_thread[(199*4)+3] <= 1'b0;
                  spc199_inst_done         <= 0;
                  spc199_phy_pc_w          <= 0;
                end else begin
                  active_thread[(199*4)]   <= 1'b1;
                  active_thread[(199*4)+1] <= 1'b1;
                  active_thread[(199*4)+2] <= 1'b1;
                  active_thread[(199*4)+3] <= 1'b1;
                  spc199_inst_done         <= `TILE199.piton_pc_vld;
                  spc199_phy_pc_w          <= `TILE199.piton_pc;
                end
            end
    

            assign spc200_thread_id = 2'b00;
            assign spc200_rtl_pc = spc200_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(200*4)]   <= 1'b0;
                  active_thread[(200*4)+1] <= 1'b0;
                  active_thread[(200*4)+2] <= 1'b0;
                  active_thread[(200*4)+3] <= 1'b0;
                  spc200_inst_done         <= 0;
                  spc200_phy_pc_w          <= 0;
                end else begin
                  active_thread[(200*4)]   <= 1'b1;
                  active_thread[(200*4)+1] <= 1'b1;
                  active_thread[(200*4)+2] <= 1'b1;
                  active_thread[(200*4)+3] <= 1'b1;
                  spc200_inst_done         <= `TILE200.piton_pc_vld;
                  spc200_phy_pc_w          <= `TILE200.piton_pc;
                end
            end
    

            assign spc201_thread_id = 2'b00;
            assign spc201_rtl_pc = spc201_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(201*4)]   <= 1'b0;
                  active_thread[(201*4)+1] <= 1'b0;
                  active_thread[(201*4)+2] <= 1'b0;
                  active_thread[(201*4)+3] <= 1'b0;
                  spc201_inst_done         <= 0;
                  spc201_phy_pc_w          <= 0;
                end else begin
                  active_thread[(201*4)]   <= 1'b1;
                  active_thread[(201*4)+1] <= 1'b1;
                  active_thread[(201*4)+2] <= 1'b1;
                  active_thread[(201*4)+3] <= 1'b1;
                  spc201_inst_done         <= `TILE201.piton_pc_vld;
                  spc201_phy_pc_w          <= `TILE201.piton_pc;
                end
            end
    

            assign spc202_thread_id = 2'b00;
            assign spc202_rtl_pc = spc202_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(202*4)]   <= 1'b0;
                  active_thread[(202*4)+1] <= 1'b0;
                  active_thread[(202*4)+2] <= 1'b0;
                  active_thread[(202*4)+3] <= 1'b0;
                  spc202_inst_done         <= 0;
                  spc202_phy_pc_w          <= 0;
                end else begin
                  active_thread[(202*4)]   <= 1'b1;
                  active_thread[(202*4)+1] <= 1'b1;
                  active_thread[(202*4)+2] <= 1'b1;
                  active_thread[(202*4)+3] <= 1'b1;
                  spc202_inst_done         <= `TILE202.piton_pc_vld;
                  spc202_phy_pc_w          <= `TILE202.piton_pc;
                end
            end
    

            assign spc203_thread_id = 2'b00;
            assign spc203_rtl_pc = spc203_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(203*4)]   <= 1'b0;
                  active_thread[(203*4)+1] <= 1'b0;
                  active_thread[(203*4)+2] <= 1'b0;
                  active_thread[(203*4)+3] <= 1'b0;
                  spc203_inst_done         <= 0;
                  spc203_phy_pc_w          <= 0;
                end else begin
                  active_thread[(203*4)]   <= 1'b1;
                  active_thread[(203*4)+1] <= 1'b1;
                  active_thread[(203*4)+2] <= 1'b1;
                  active_thread[(203*4)+3] <= 1'b1;
                  spc203_inst_done         <= `TILE203.piton_pc_vld;
                  spc203_phy_pc_w          <= `TILE203.piton_pc;
                end
            end
    

            assign spc204_thread_id = 2'b00;
            assign spc204_rtl_pc = spc204_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(204*4)]   <= 1'b0;
                  active_thread[(204*4)+1] <= 1'b0;
                  active_thread[(204*4)+2] <= 1'b0;
                  active_thread[(204*4)+3] <= 1'b0;
                  spc204_inst_done         <= 0;
                  spc204_phy_pc_w          <= 0;
                end else begin
                  active_thread[(204*4)]   <= 1'b1;
                  active_thread[(204*4)+1] <= 1'b1;
                  active_thread[(204*4)+2] <= 1'b1;
                  active_thread[(204*4)+3] <= 1'b1;
                  spc204_inst_done         <= `TILE204.piton_pc_vld;
                  spc204_phy_pc_w          <= `TILE204.piton_pc;
                end
            end
    

            assign spc205_thread_id = 2'b00;
            assign spc205_rtl_pc = spc205_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(205*4)]   <= 1'b0;
                  active_thread[(205*4)+1] <= 1'b0;
                  active_thread[(205*4)+2] <= 1'b0;
                  active_thread[(205*4)+3] <= 1'b0;
                  spc205_inst_done         <= 0;
                  spc205_phy_pc_w          <= 0;
                end else begin
                  active_thread[(205*4)]   <= 1'b1;
                  active_thread[(205*4)+1] <= 1'b1;
                  active_thread[(205*4)+2] <= 1'b1;
                  active_thread[(205*4)+3] <= 1'b1;
                  spc205_inst_done         <= `TILE205.piton_pc_vld;
                  spc205_phy_pc_w          <= `TILE205.piton_pc;
                end
            end
    

            assign spc206_thread_id = 2'b00;
            assign spc206_rtl_pc = spc206_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(206*4)]   <= 1'b0;
                  active_thread[(206*4)+1] <= 1'b0;
                  active_thread[(206*4)+2] <= 1'b0;
                  active_thread[(206*4)+3] <= 1'b0;
                  spc206_inst_done         <= 0;
                  spc206_phy_pc_w          <= 0;
                end else begin
                  active_thread[(206*4)]   <= 1'b1;
                  active_thread[(206*4)+1] <= 1'b1;
                  active_thread[(206*4)+2] <= 1'b1;
                  active_thread[(206*4)+3] <= 1'b1;
                  spc206_inst_done         <= `TILE206.piton_pc_vld;
                  spc206_phy_pc_w          <= `TILE206.piton_pc;
                end
            end
    

            assign spc207_thread_id = 2'b00;
            assign spc207_rtl_pc = spc207_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(207*4)]   <= 1'b0;
                  active_thread[(207*4)+1] <= 1'b0;
                  active_thread[(207*4)+2] <= 1'b0;
                  active_thread[(207*4)+3] <= 1'b0;
                  spc207_inst_done         <= 0;
                  spc207_phy_pc_w          <= 0;
                end else begin
                  active_thread[(207*4)]   <= 1'b1;
                  active_thread[(207*4)+1] <= 1'b1;
                  active_thread[(207*4)+2] <= 1'b1;
                  active_thread[(207*4)+3] <= 1'b1;
                  spc207_inst_done         <= `TILE207.piton_pc_vld;
                  spc207_phy_pc_w          <= `TILE207.piton_pc;
                end
            end
    

            assign spc208_thread_id = 2'b00;
            assign spc208_rtl_pc = spc208_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(208*4)]   <= 1'b0;
                  active_thread[(208*4)+1] <= 1'b0;
                  active_thread[(208*4)+2] <= 1'b0;
                  active_thread[(208*4)+3] <= 1'b0;
                  spc208_inst_done         <= 0;
                  spc208_phy_pc_w          <= 0;
                end else begin
                  active_thread[(208*4)]   <= 1'b1;
                  active_thread[(208*4)+1] <= 1'b1;
                  active_thread[(208*4)+2] <= 1'b1;
                  active_thread[(208*4)+3] <= 1'b1;
                  spc208_inst_done         <= `TILE208.piton_pc_vld;
                  spc208_phy_pc_w          <= `TILE208.piton_pc;
                end
            end
    

            assign spc209_thread_id = 2'b00;
            assign spc209_rtl_pc = spc209_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(209*4)]   <= 1'b0;
                  active_thread[(209*4)+1] <= 1'b0;
                  active_thread[(209*4)+2] <= 1'b0;
                  active_thread[(209*4)+3] <= 1'b0;
                  spc209_inst_done         <= 0;
                  spc209_phy_pc_w          <= 0;
                end else begin
                  active_thread[(209*4)]   <= 1'b1;
                  active_thread[(209*4)+1] <= 1'b1;
                  active_thread[(209*4)+2] <= 1'b1;
                  active_thread[(209*4)+3] <= 1'b1;
                  spc209_inst_done         <= `TILE209.piton_pc_vld;
                  spc209_phy_pc_w          <= `TILE209.piton_pc;
                end
            end
    

            assign spc210_thread_id = 2'b00;
            assign spc210_rtl_pc = spc210_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(210*4)]   <= 1'b0;
                  active_thread[(210*4)+1] <= 1'b0;
                  active_thread[(210*4)+2] <= 1'b0;
                  active_thread[(210*4)+3] <= 1'b0;
                  spc210_inst_done         <= 0;
                  spc210_phy_pc_w          <= 0;
                end else begin
                  active_thread[(210*4)]   <= 1'b1;
                  active_thread[(210*4)+1] <= 1'b1;
                  active_thread[(210*4)+2] <= 1'b1;
                  active_thread[(210*4)+3] <= 1'b1;
                  spc210_inst_done         <= `TILE210.piton_pc_vld;
                  spc210_phy_pc_w          <= `TILE210.piton_pc;
                end
            end
    

            assign spc211_thread_id = 2'b00;
            assign spc211_rtl_pc = spc211_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(211*4)]   <= 1'b0;
                  active_thread[(211*4)+1] <= 1'b0;
                  active_thread[(211*4)+2] <= 1'b0;
                  active_thread[(211*4)+3] <= 1'b0;
                  spc211_inst_done         <= 0;
                  spc211_phy_pc_w          <= 0;
                end else begin
                  active_thread[(211*4)]   <= 1'b1;
                  active_thread[(211*4)+1] <= 1'b1;
                  active_thread[(211*4)+2] <= 1'b1;
                  active_thread[(211*4)+3] <= 1'b1;
                  spc211_inst_done         <= `TILE211.piton_pc_vld;
                  spc211_phy_pc_w          <= `TILE211.piton_pc;
                end
            end
    

            assign spc212_thread_id = 2'b00;
            assign spc212_rtl_pc = spc212_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(212*4)]   <= 1'b0;
                  active_thread[(212*4)+1] <= 1'b0;
                  active_thread[(212*4)+2] <= 1'b0;
                  active_thread[(212*4)+3] <= 1'b0;
                  spc212_inst_done         <= 0;
                  spc212_phy_pc_w          <= 0;
                end else begin
                  active_thread[(212*4)]   <= 1'b1;
                  active_thread[(212*4)+1] <= 1'b1;
                  active_thread[(212*4)+2] <= 1'b1;
                  active_thread[(212*4)+3] <= 1'b1;
                  spc212_inst_done         <= `TILE212.piton_pc_vld;
                  spc212_phy_pc_w          <= `TILE212.piton_pc;
                end
            end
    

            assign spc213_thread_id = 2'b00;
            assign spc213_rtl_pc = spc213_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(213*4)]   <= 1'b0;
                  active_thread[(213*4)+1] <= 1'b0;
                  active_thread[(213*4)+2] <= 1'b0;
                  active_thread[(213*4)+3] <= 1'b0;
                  spc213_inst_done         <= 0;
                  spc213_phy_pc_w          <= 0;
                end else begin
                  active_thread[(213*4)]   <= 1'b1;
                  active_thread[(213*4)+1] <= 1'b1;
                  active_thread[(213*4)+2] <= 1'b1;
                  active_thread[(213*4)+3] <= 1'b1;
                  spc213_inst_done         <= `TILE213.piton_pc_vld;
                  spc213_phy_pc_w          <= `TILE213.piton_pc;
                end
            end
    

            assign spc214_thread_id = 2'b00;
            assign spc214_rtl_pc = spc214_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(214*4)]   <= 1'b0;
                  active_thread[(214*4)+1] <= 1'b0;
                  active_thread[(214*4)+2] <= 1'b0;
                  active_thread[(214*4)+3] <= 1'b0;
                  spc214_inst_done         <= 0;
                  spc214_phy_pc_w          <= 0;
                end else begin
                  active_thread[(214*4)]   <= 1'b1;
                  active_thread[(214*4)+1] <= 1'b1;
                  active_thread[(214*4)+2] <= 1'b1;
                  active_thread[(214*4)+3] <= 1'b1;
                  spc214_inst_done         <= `TILE214.piton_pc_vld;
                  spc214_phy_pc_w          <= `TILE214.piton_pc;
                end
            end
    

            assign spc215_thread_id = 2'b00;
            assign spc215_rtl_pc = spc215_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(215*4)]   <= 1'b0;
                  active_thread[(215*4)+1] <= 1'b0;
                  active_thread[(215*4)+2] <= 1'b0;
                  active_thread[(215*4)+3] <= 1'b0;
                  spc215_inst_done         <= 0;
                  spc215_phy_pc_w          <= 0;
                end else begin
                  active_thread[(215*4)]   <= 1'b1;
                  active_thread[(215*4)+1] <= 1'b1;
                  active_thread[(215*4)+2] <= 1'b1;
                  active_thread[(215*4)+3] <= 1'b1;
                  spc215_inst_done         <= `TILE215.piton_pc_vld;
                  spc215_phy_pc_w          <= `TILE215.piton_pc;
                end
            end
    

            assign spc216_thread_id = 2'b00;
            assign spc216_rtl_pc = spc216_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(216*4)]   <= 1'b0;
                  active_thread[(216*4)+1] <= 1'b0;
                  active_thread[(216*4)+2] <= 1'b0;
                  active_thread[(216*4)+3] <= 1'b0;
                  spc216_inst_done         <= 0;
                  spc216_phy_pc_w          <= 0;
                end else begin
                  active_thread[(216*4)]   <= 1'b1;
                  active_thread[(216*4)+1] <= 1'b1;
                  active_thread[(216*4)+2] <= 1'b1;
                  active_thread[(216*4)+3] <= 1'b1;
                  spc216_inst_done         <= `TILE216.piton_pc_vld;
                  spc216_phy_pc_w          <= `TILE216.piton_pc;
                end
            end
    

            assign spc217_thread_id = 2'b00;
            assign spc217_rtl_pc = spc217_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(217*4)]   <= 1'b0;
                  active_thread[(217*4)+1] <= 1'b0;
                  active_thread[(217*4)+2] <= 1'b0;
                  active_thread[(217*4)+3] <= 1'b0;
                  spc217_inst_done         <= 0;
                  spc217_phy_pc_w          <= 0;
                end else begin
                  active_thread[(217*4)]   <= 1'b1;
                  active_thread[(217*4)+1] <= 1'b1;
                  active_thread[(217*4)+2] <= 1'b1;
                  active_thread[(217*4)+3] <= 1'b1;
                  spc217_inst_done         <= `TILE217.piton_pc_vld;
                  spc217_phy_pc_w          <= `TILE217.piton_pc;
                end
            end
    

            assign spc218_thread_id = 2'b00;
            assign spc218_rtl_pc = spc218_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(218*4)]   <= 1'b0;
                  active_thread[(218*4)+1] <= 1'b0;
                  active_thread[(218*4)+2] <= 1'b0;
                  active_thread[(218*4)+3] <= 1'b0;
                  spc218_inst_done         <= 0;
                  spc218_phy_pc_w          <= 0;
                end else begin
                  active_thread[(218*4)]   <= 1'b1;
                  active_thread[(218*4)+1] <= 1'b1;
                  active_thread[(218*4)+2] <= 1'b1;
                  active_thread[(218*4)+3] <= 1'b1;
                  spc218_inst_done         <= `TILE218.piton_pc_vld;
                  spc218_phy_pc_w          <= `TILE218.piton_pc;
                end
            end
    

            assign spc219_thread_id = 2'b00;
            assign spc219_rtl_pc = spc219_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(219*4)]   <= 1'b0;
                  active_thread[(219*4)+1] <= 1'b0;
                  active_thread[(219*4)+2] <= 1'b0;
                  active_thread[(219*4)+3] <= 1'b0;
                  spc219_inst_done         <= 0;
                  spc219_phy_pc_w          <= 0;
                end else begin
                  active_thread[(219*4)]   <= 1'b1;
                  active_thread[(219*4)+1] <= 1'b1;
                  active_thread[(219*4)+2] <= 1'b1;
                  active_thread[(219*4)+3] <= 1'b1;
                  spc219_inst_done         <= `TILE219.piton_pc_vld;
                  spc219_phy_pc_w          <= `TILE219.piton_pc;
                end
            end
    

            assign spc220_thread_id = 2'b00;
            assign spc220_rtl_pc = spc220_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(220*4)]   <= 1'b0;
                  active_thread[(220*4)+1] <= 1'b0;
                  active_thread[(220*4)+2] <= 1'b0;
                  active_thread[(220*4)+3] <= 1'b0;
                  spc220_inst_done         <= 0;
                  spc220_phy_pc_w          <= 0;
                end else begin
                  active_thread[(220*4)]   <= 1'b1;
                  active_thread[(220*4)+1] <= 1'b1;
                  active_thread[(220*4)+2] <= 1'b1;
                  active_thread[(220*4)+3] <= 1'b1;
                  spc220_inst_done         <= `TILE220.piton_pc_vld;
                  spc220_phy_pc_w          <= `TILE220.piton_pc;
                end
            end
    

            assign spc221_thread_id = 2'b00;
            assign spc221_rtl_pc = spc221_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(221*4)]   <= 1'b0;
                  active_thread[(221*4)+1] <= 1'b0;
                  active_thread[(221*4)+2] <= 1'b0;
                  active_thread[(221*4)+3] <= 1'b0;
                  spc221_inst_done         <= 0;
                  spc221_phy_pc_w          <= 0;
                end else begin
                  active_thread[(221*4)]   <= 1'b1;
                  active_thread[(221*4)+1] <= 1'b1;
                  active_thread[(221*4)+2] <= 1'b1;
                  active_thread[(221*4)+3] <= 1'b1;
                  spc221_inst_done         <= `TILE221.piton_pc_vld;
                  spc221_phy_pc_w          <= `TILE221.piton_pc;
                end
            end
    

            assign spc222_thread_id = 2'b00;
            assign spc222_rtl_pc = spc222_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(222*4)]   <= 1'b0;
                  active_thread[(222*4)+1] <= 1'b0;
                  active_thread[(222*4)+2] <= 1'b0;
                  active_thread[(222*4)+3] <= 1'b0;
                  spc222_inst_done         <= 0;
                  spc222_phy_pc_w          <= 0;
                end else begin
                  active_thread[(222*4)]   <= 1'b1;
                  active_thread[(222*4)+1] <= 1'b1;
                  active_thread[(222*4)+2] <= 1'b1;
                  active_thread[(222*4)+3] <= 1'b1;
                  spc222_inst_done         <= `TILE222.piton_pc_vld;
                  spc222_phy_pc_w          <= `TILE222.piton_pc;
                end
            end
    

            assign spc223_thread_id = 2'b00;
            assign spc223_rtl_pc = spc223_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(223*4)]   <= 1'b0;
                  active_thread[(223*4)+1] <= 1'b0;
                  active_thread[(223*4)+2] <= 1'b0;
                  active_thread[(223*4)+3] <= 1'b0;
                  spc223_inst_done         <= 0;
                  spc223_phy_pc_w          <= 0;
                end else begin
                  active_thread[(223*4)]   <= 1'b1;
                  active_thread[(223*4)+1] <= 1'b1;
                  active_thread[(223*4)+2] <= 1'b1;
                  active_thread[(223*4)+3] <= 1'b1;
                  spc223_inst_done         <= `TILE223.piton_pc_vld;
                  spc223_phy_pc_w          <= `TILE223.piton_pc;
                end
            end
    

            assign spc224_thread_id = 2'b00;
            assign spc224_rtl_pc = spc224_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(224*4)]   <= 1'b0;
                  active_thread[(224*4)+1] <= 1'b0;
                  active_thread[(224*4)+2] <= 1'b0;
                  active_thread[(224*4)+3] <= 1'b0;
                  spc224_inst_done         <= 0;
                  spc224_phy_pc_w          <= 0;
                end else begin
                  active_thread[(224*4)]   <= 1'b1;
                  active_thread[(224*4)+1] <= 1'b1;
                  active_thread[(224*4)+2] <= 1'b1;
                  active_thread[(224*4)+3] <= 1'b1;
                  spc224_inst_done         <= `TILE224.piton_pc_vld;
                  spc224_phy_pc_w          <= `TILE224.piton_pc;
                end
            end
    

            assign spc225_thread_id = 2'b00;
            assign spc225_rtl_pc = spc225_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(225*4)]   <= 1'b0;
                  active_thread[(225*4)+1] <= 1'b0;
                  active_thread[(225*4)+2] <= 1'b0;
                  active_thread[(225*4)+3] <= 1'b0;
                  spc225_inst_done         <= 0;
                  spc225_phy_pc_w          <= 0;
                end else begin
                  active_thread[(225*4)]   <= 1'b1;
                  active_thread[(225*4)+1] <= 1'b1;
                  active_thread[(225*4)+2] <= 1'b1;
                  active_thread[(225*4)+3] <= 1'b1;
                  spc225_inst_done         <= `TILE225.piton_pc_vld;
                  spc225_phy_pc_w          <= `TILE225.piton_pc;
                end
            end
    

            assign spc226_thread_id = 2'b00;
            assign spc226_rtl_pc = spc226_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(226*4)]   <= 1'b0;
                  active_thread[(226*4)+1] <= 1'b0;
                  active_thread[(226*4)+2] <= 1'b0;
                  active_thread[(226*4)+3] <= 1'b0;
                  spc226_inst_done         <= 0;
                  spc226_phy_pc_w          <= 0;
                end else begin
                  active_thread[(226*4)]   <= 1'b1;
                  active_thread[(226*4)+1] <= 1'b1;
                  active_thread[(226*4)+2] <= 1'b1;
                  active_thread[(226*4)+3] <= 1'b1;
                  spc226_inst_done         <= `TILE226.piton_pc_vld;
                  spc226_phy_pc_w          <= `TILE226.piton_pc;
                end
            end
    

            assign spc227_thread_id = 2'b00;
            assign spc227_rtl_pc = spc227_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(227*4)]   <= 1'b0;
                  active_thread[(227*4)+1] <= 1'b0;
                  active_thread[(227*4)+2] <= 1'b0;
                  active_thread[(227*4)+3] <= 1'b0;
                  spc227_inst_done         <= 0;
                  spc227_phy_pc_w          <= 0;
                end else begin
                  active_thread[(227*4)]   <= 1'b1;
                  active_thread[(227*4)+1] <= 1'b1;
                  active_thread[(227*4)+2] <= 1'b1;
                  active_thread[(227*4)+3] <= 1'b1;
                  spc227_inst_done         <= `TILE227.piton_pc_vld;
                  spc227_phy_pc_w          <= `TILE227.piton_pc;
                end
            end
    

            assign spc228_thread_id = 2'b00;
            assign spc228_rtl_pc = spc228_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(228*4)]   <= 1'b0;
                  active_thread[(228*4)+1] <= 1'b0;
                  active_thread[(228*4)+2] <= 1'b0;
                  active_thread[(228*4)+3] <= 1'b0;
                  spc228_inst_done         <= 0;
                  spc228_phy_pc_w          <= 0;
                end else begin
                  active_thread[(228*4)]   <= 1'b1;
                  active_thread[(228*4)+1] <= 1'b1;
                  active_thread[(228*4)+2] <= 1'b1;
                  active_thread[(228*4)+3] <= 1'b1;
                  spc228_inst_done         <= `TILE228.piton_pc_vld;
                  spc228_phy_pc_w          <= `TILE228.piton_pc;
                end
            end
    

            assign spc229_thread_id = 2'b00;
            assign spc229_rtl_pc = spc229_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(229*4)]   <= 1'b0;
                  active_thread[(229*4)+1] <= 1'b0;
                  active_thread[(229*4)+2] <= 1'b0;
                  active_thread[(229*4)+3] <= 1'b0;
                  spc229_inst_done         <= 0;
                  spc229_phy_pc_w          <= 0;
                end else begin
                  active_thread[(229*4)]   <= 1'b1;
                  active_thread[(229*4)+1] <= 1'b1;
                  active_thread[(229*4)+2] <= 1'b1;
                  active_thread[(229*4)+3] <= 1'b1;
                  spc229_inst_done         <= `TILE229.piton_pc_vld;
                  spc229_phy_pc_w          <= `TILE229.piton_pc;
                end
            end
    

            assign spc230_thread_id = 2'b00;
            assign spc230_rtl_pc = spc230_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(230*4)]   <= 1'b0;
                  active_thread[(230*4)+1] <= 1'b0;
                  active_thread[(230*4)+2] <= 1'b0;
                  active_thread[(230*4)+3] <= 1'b0;
                  spc230_inst_done         <= 0;
                  spc230_phy_pc_w          <= 0;
                end else begin
                  active_thread[(230*4)]   <= 1'b1;
                  active_thread[(230*4)+1] <= 1'b1;
                  active_thread[(230*4)+2] <= 1'b1;
                  active_thread[(230*4)+3] <= 1'b1;
                  spc230_inst_done         <= `TILE230.piton_pc_vld;
                  spc230_phy_pc_w          <= `TILE230.piton_pc;
                end
            end
    

            assign spc231_thread_id = 2'b00;
            assign spc231_rtl_pc = spc231_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(231*4)]   <= 1'b0;
                  active_thread[(231*4)+1] <= 1'b0;
                  active_thread[(231*4)+2] <= 1'b0;
                  active_thread[(231*4)+3] <= 1'b0;
                  spc231_inst_done         <= 0;
                  spc231_phy_pc_w          <= 0;
                end else begin
                  active_thread[(231*4)]   <= 1'b1;
                  active_thread[(231*4)+1] <= 1'b1;
                  active_thread[(231*4)+2] <= 1'b1;
                  active_thread[(231*4)+3] <= 1'b1;
                  spc231_inst_done         <= `TILE231.piton_pc_vld;
                  spc231_phy_pc_w          <= `TILE231.piton_pc;
                end
            end
    

            assign spc232_thread_id = 2'b00;
            assign spc232_rtl_pc = spc232_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(232*4)]   <= 1'b0;
                  active_thread[(232*4)+1] <= 1'b0;
                  active_thread[(232*4)+2] <= 1'b0;
                  active_thread[(232*4)+3] <= 1'b0;
                  spc232_inst_done         <= 0;
                  spc232_phy_pc_w          <= 0;
                end else begin
                  active_thread[(232*4)]   <= 1'b1;
                  active_thread[(232*4)+1] <= 1'b1;
                  active_thread[(232*4)+2] <= 1'b1;
                  active_thread[(232*4)+3] <= 1'b1;
                  spc232_inst_done         <= `TILE232.piton_pc_vld;
                  spc232_phy_pc_w          <= `TILE232.piton_pc;
                end
            end
    

            assign spc233_thread_id = 2'b00;
            assign spc233_rtl_pc = spc233_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(233*4)]   <= 1'b0;
                  active_thread[(233*4)+1] <= 1'b0;
                  active_thread[(233*4)+2] <= 1'b0;
                  active_thread[(233*4)+3] <= 1'b0;
                  spc233_inst_done         <= 0;
                  spc233_phy_pc_w          <= 0;
                end else begin
                  active_thread[(233*4)]   <= 1'b1;
                  active_thread[(233*4)+1] <= 1'b1;
                  active_thread[(233*4)+2] <= 1'b1;
                  active_thread[(233*4)+3] <= 1'b1;
                  spc233_inst_done         <= `TILE233.piton_pc_vld;
                  spc233_phy_pc_w          <= `TILE233.piton_pc;
                end
            end
    

            assign spc234_thread_id = 2'b00;
            assign spc234_rtl_pc = spc234_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(234*4)]   <= 1'b0;
                  active_thread[(234*4)+1] <= 1'b0;
                  active_thread[(234*4)+2] <= 1'b0;
                  active_thread[(234*4)+3] <= 1'b0;
                  spc234_inst_done         <= 0;
                  spc234_phy_pc_w          <= 0;
                end else begin
                  active_thread[(234*4)]   <= 1'b1;
                  active_thread[(234*4)+1] <= 1'b1;
                  active_thread[(234*4)+2] <= 1'b1;
                  active_thread[(234*4)+3] <= 1'b1;
                  spc234_inst_done         <= `TILE234.piton_pc_vld;
                  spc234_phy_pc_w          <= `TILE234.piton_pc;
                end
            end
    

            assign spc235_thread_id = 2'b00;
            assign spc235_rtl_pc = spc235_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(235*4)]   <= 1'b0;
                  active_thread[(235*4)+1] <= 1'b0;
                  active_thread[(235*4)+2] <= 1'b0;
                  active_thread[(235*4)+3] <= 1'b0;
                  spc235_inst_done         <= 0;
                  spc235_phy_pc_w          <= 0;
                end else begin
                  active_thread[(235*4)]   <= 1'b1;
                  active_thread[(235*4)+1] <= 1'b1;
                  active_thread[(235*4)+2] <= 1'b1;
                  active_thread[(235*4)+3] <= 1'b1;
                  spc235_inst_done         <= `TILE235.piton_pc_vld;
                  spc235_phy_pc_w          <= `TILE235.piton_pc;
                end
            end
    

            assign spc236_thread_id = 2'b00;
            assign spc236_rtl_pc = spc236_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(236*4)]   <= 1'b0;
                  active_thread[(236*4)+1] <= 1'b0;
                  active_thread[(236*4)+2] <= 1'b0;
                  active_thread[(236*4)+3] <= 1'b0;
                  spc236_inst_done         <= 0;
                  spc236_phy_pc_w          <= 0;
                end else begin
                  active_thread[(236*4)]   <= 1'b1;
                  active_thread[(236*4)+1] <= 1'b1;
                  active_thread[(236*4)+2] <= 1'b1;
                  active_thread[(236*4)+3] <= 1'b1;
                  spc236_inst_done         <= `TILE236.piton_pc_vld;
                  spc236_phy_pc_w          <= `TILE236.piton_pc;
                end
            end
    

            assign spc237_thread_id = 2'b00;
            assign spc237_rtl_pc = spc237_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(237*4)]   <= 1'b0;
                  active_thread[(237*4)+1] <= 1'b0;
                  active_thread[(237*4)+2] <= 1'b0;
                  active_thread[(237*4)+3] <= 1'b0;
                  spc237_inst_done         <= 0;
                  spc237_phy_pc_w          <= 0;
                end else begin
                  active_thread[(237*4)]   <= 1'b1;
                  active_thread[(237*4)+1] <= 1'b1;
                  active_thread[(237*4)+2] <= 1'b1;
                  active_thread[(237*4)+3] <= 1'b1;
                  spc237_inst_done         <= `TILE237.piton_pc_vld;
                  spc237_phy_pc_w          <= `TILE237.piton_pc;
                end
            end
    

            assign spc238_thread_id = 2'b00;
            assign spc238_rtl_pc = spc238_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(238*4)]   <= 1'b0;
                  active_thread[(238*4)+1] <= 1'b0;
                  active_thread[(238*4)+2] <= 1'b0;
                  active_thread[(238*4)+3] <= 1'b0;
                  spc238_inst_done         <= 0;
                  spc238_phy_pc_w          <= 0;
                end else begin
                  active_thread[(238*4)]   <= 1'b1;
                  active_thread[(238*4)+1] <= 1'b1;
                  active_thread[(238*4)+2] <= 1'b1;
                  active_thread[(238*4)+3] <= 1'b1;
                  spc238_inst_done         <= `TILE238.piton_pc_vld;
                  spc238_phy_pc_w          <= `TILE238.piton_pc;
                end
            end
    

            assign spc239_thread_id = 2'b00;
            assign spc239_rtl_pc = spc239_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(239*4)]   <= 1'b0;
                  active_thread[(239*4)+1] <= 1'b0;
                  active_thread[(239*4)+2] <= 1'b0;
                  active_thread[(239*4)+3] <= 1'b0;
                  spc239_inst_done         <= 0;
                  spc239_phy_pc_w          <= 0;
                end else begin
                  active_thread[(239*4)]   <= 1'b1;
                  active_thread[(239*4)+1] <= 1'b1;
                  active_thread[(239*4)+2] <= 1'b1;
                  active_thread[(239*4)+3] <= 1'b1;
                  spc239_inst_done         <= `TILE239.piton_pc_vld;
                  spc239_phy_pc_w          <= `TILE239.piton_pc;
                end
            end
    

            assign spc240_thread_id = 2'b00;
            assign spc240_rtl_pc = spc240_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(240*4)]   <= 1'b0;
                  active_thread[(240*4)+1] <= 1'b0;
                  active_thread[(240*4)+2] <= 1'b0;
                  active_thread[(240*4)+3] <= 1'b0;
                  spc240_inst_done         <= 0;
                  spc240_phy_pc_w          <= 0;
                end else begin
                  active_thread[(240*4)]   <= 1'b1;
                  active_thread[(240*4)+1] <= 1'b1;
                  active_thread[(240*4)+2] <= 1'b1;
                  active_thread[(240*4)+3] <= 1'b1;
                  spc240_inst_done         <= `TILE240.piton_pc_vld;
                  spc240_phy_pc_w          <= `TILE240.piton_pc;
                end
            end
    

            assign spc241_thread_id = 2'b00;
            assign spc241_rtl_pc = spc241_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(241*4)]   <= 1'b0;
                  active_thread[(241*4)+1] <= 1'b0;
                  active_thread[(241*4)+2] <= 1'b0;
                  active_thread[(241*4)+3] <= 1'b0;
                  spc241_inst_done         <= 0;
                  spc241_phy_pc_w          <= 0;
                end else begin
                  active_thread[(241*4)]   <= 1'b1;
                  active_thread[(241*4)+1] <= 1'b1;
                  active_thread[(241*4)+2] <= 1'b1;
                  active_thread[(241*4)+3] <= 1'b1;
                  spc241_inst_done         <= `TILE241.piton_pc_vld;
                  spc241_phy_pc_w          <= `TILE241.piton_pc;
                end
            end
    

            assign spc242_thread_id = 2'b00;
            assign spc242_rtl_pc = spc242_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(242*4)]   <= 1'b0;
                  active_thread[(242*4)+1] <= 1'b0;
                  active_thread[(242*4)+2] <= 1'b0;
                  active_thread[(242*4)+3] <= 1'b0;
                  spc242_inst_done         <= 0;
                  spc242_phy_pc_w          <= 0;
                end else begin
                  active_thread[(242*4)]   <= 1'b1;
                  active_thread[(242*4)+1] <= 1'b1;
                  active_thread[(242*4)+2] <= 1'b1;
                  active_thread[(242*4)+3] <= 1'b1;
                  spc242_inst_done         <= `TILE242.piton_pc_vld;
                  spc242_phy_pc_w          <= `TILE242.piton_pc;
                end
            end
    

            assign spc243_thread_id = 2'b00;
            assign spc243_rtl_pc = spc243_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(243*4)]   <= 1'b0;
                  active_thread[(243*4)+1] <= 1'b0;
                  active_thread[(243*4)+2] <= 1'b0;
                  active_thread[(243*4)+3] <= 1'b0;
                  spc243_inst_done         <= 0;
                  spc243_phy_pc_w          <= 0;
                end else begin
                  active_thread[(243*4)]   <= 1'b1;
                  active_thread[(243*4)+1] <= 1'b1;
                  active_thread[(243*4)+2] <= 1'b1;
                  active_thread[(243*4)+3] <= 1'b1;
                  spc243_inst_done         <= `TILE243.piton_pc_vld;
                  spc243_phy_pc_w          <= `TILE243.piton_pc;
                end
            end
    

            assign spc244_thread_id = 2'b00;
            assign spc244_rtl_pc = spc244_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(244*4)]   <= 1'b0;
                  active_thread[(244*4)+1] <= 1'b0;
                  active_thread[(244*4)+2] <= 1'b0;
                  active_thread[(244*4)+3] <= 1'b0;
                  spc244_inst_done         <= 0;
                  spc244_phy_pc_w          <= 0;
                end else begin
                  active_thread[(244*4)]   <= 1'b1;
                  active_thread[(244*4)+1] <= 1'b1;
                  active_thread[(244*4)+2] <= 1'b1;
                  active_thread[(244*4)+3] <= 1'b1;
                  spc244_inst_done         <= `TILE244.piton_pc_vld;
                  spc244_phy_pc_w          <= `TILE244.piton_pc;
                end
            end
    

            assign spc245_thread_id = 2'b00;
            assign spc245_rtl_pc = spc245_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(245*4)]   <= 1'b0;
                  active_thread[(245*4)+1] <= 1'b0;
                  active_thread[(245*4)+2] <= 1'b0;
                  active_thread[(245*4)+3] <= 1'b0;
                  spc245_inst_done         <= 0;
                  spc245_phy_pc_w          <= 0;
                end else begin
                  active_thread[(245*4)]   <= 1'b1;
                  active_thread[(245*4)+1] <= 1'b1;
                  active_thread[(245*4)+2] <= 1'b1;
                  active_thread[(245*4)+3] <= 1'b1;
                  spc245_inst_done         <= `TILE245.piton_pc_vld;
                  spc245_phy_pc_w          <= `TILE245.piton_pc;
                end
            end
    

            assign spc246_thread_id = 2'b00;
            assign spc246_rtl_pc = spc246_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(246*4)]   <= 1'b0;
                  active_thread[(246*4)+1] <= 1'b0;
                  active_thread[(246*4)+2] <= 1'b0;
                  active_thread[(246*4)+3] <= 1'b0;
                  spc246_inst_done         <= 0;
                  spc246_phy_pc_w          <= 0;
                end else begin
                  active_thread[(246*4)]   <= 1'b1;
                  active_thread[(246*4)+1] <= 1'b1;
                  active_thread[(246*4)+2] <= 1'b1;
                  active_thread[(246*4)+3] <= 1'b1;
                  spc246_inst_done         <= `TILE246.piton_pc_vld;
                  spc246_phy_pc_w          <= `TILE246.piton_pc;
                end
            end
    

            assign spc247_thread_id = 2'b00;
            assign spc247_rtl_pc = spc247_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(247*4)]   <= 1'b0;
                  active_thread[(247*4)+1] <= 1'b0;
                  active_thread[(247*4)+2] <= 1'b0;
                  active_thread[(247*4)+3] <= 1'b0;
                  spc247_inst_done         <= 0;
                  spc247_phy_pc_w          <= 0;
                end else begin
                  active_thread[(247*4)]   <= 1'b1;
                  active_thread[(247*4)+1] <= 1'b1;
                  active_thread[(247*4)+2] <= 1'b1;
                  active_thread[(247*4)+3] <= 1'b1;
                  spc247_inst_done         <= `TILE247.piton_pc_vld;
                  spc247_phy_pc_w          <= `TILE247.piton_pc;
                end
            end
    

            assign spc248_thread_id = 2'b00;
            assign spc248_rtl_pc = spc248_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(248*4)]   <= 1'b0;
                  active_thread[(248*4)+1] <= 1'b0;
                  active_thread[(248*4)+2] <= 1'b0;
                  active_thread[(248*4)+3] <= 1'b0;
                  spc248_inst_done         <= 0;
                  spc248_phy_pc_w          <= 0;
                end else begin
                  active_thread[(248*4)]   <= 1'b1;
                  active_thread[(248*4)+1] <= 1'b1;
                  active_thread[(248*4)+2] <= 1'b1;
                  active_thread[(248*4)+3] <= 1'b1;
                  spc248_inst_done         <= `TILE248.piton_pc_vld;
                  spc248_phy_pc_w          <= `TILE248.piton_pc;
                end
            end
    

            assign spc249_thread_id = 2'b00;
            assign spc249_rtl_pc = spc249_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(249*4)]   <= 1'b0;
                  active_thread[(249*4)+1] <= 1'b0;
                  active_thread[(249*4)+2] <= 1'b0;
                  active_thread[(249*4)+3] <= 1'b0;
                  spc249_inst_done         <= 0;
                  spc249_phy_pc_w          <= 0;
                end else begin
                  active_thread[(249*4)]   <= 1'b1;
                  active_thread[(249*4)+1] <= 1'b1;
                  active_thread[(249*4)+2] <= 1'b1;
                  active_thread[(249*4)+3] <= 1'b1;
                  spc249_inst_done         <= `TILE249.piton_pc_vld;
                  spc249_phy_pc_w          <= `TILE249.piton_pc;
                end
            end
    

            assign spc250_thread_id = 2'b00;
            assign spc250_rtl_pc = spc250_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(250*4)]   <= 1'b0;
                  active_thread[(250*4)+1] <= 1'b0;
                  active_thread[(250*4)+2] <= 1'b0;
                  active_thread[(250*4)+3] <= 1'b0;
                  spc250_inst_done         <= 0;
                  spc250_phy_pc_w          <= 0;
                end else begin
                  active_thread[(250*4)]   <= 1'b1;
                  active_thread[(250*4)+1] <= 1'b1;
                  active_thread[(250*4)+2] <= 1'b1;
                  active_thread[(250*4)+3] <= 1'b1;
                  spc250_inst_done         <= `TILE250.piton_pc_vld;
                  spc250_phy_pc_w          <= `TILE250.piton_pc;
                end
            end
    

            assign spc251_thread_id = 2'b00;
            assign spc251_rtl_pc = spc251_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(251*4)]   <= 1'b0;
                  active_thread[(251*4)+1] <= 1'b0;
                  active_thread[(251*4)+2] <= 1'b0;
                  active_thread[(251*4)+3] <= 1'b0;
                  spc251_inst_done         <= 0;
                  spc251_phy_pc_w          <= 0;
                end else begin
                  active_thread[(251*4)]   <= 1'b1;
                  active_thread[(251*4)+1] <= 1'b1;
                  active_thread[(251*4)+2] <= 1'b1;
                  active_thread[(251*4)+3] <= 1'b1;
                  spc251_inst_done         <= `TILE251.piton_pc_vld;
                  spc251_phy_pc_w          <= `TILE251.piton_pc;
                end
            end
    

            assign spc252_thread_id = 2'b00;
            assign spc252_rtl_pc = spc252_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(252*4)]   <= 1'b0;
                  active_thread[(252*4)+1] <= 1'b0;
                  active_thread[(252*4)+2] <= 1'b0;
                  active_thread[(252*4)+3] <= 1'b0;
                  spc252_inst_done         <= 0;
                  spc252_phy_pc_w          <= 0;
                end else begin
                  active_thread[(252*4)]   <= 1'b1;
                  active_thread[(252*4)+1] <= 1'b1;
                  active_thread[(252*4)+2] <= 1'b1;
                  active_thread[(252*4)+3] <= 1'b1;
                  spc252_inst_done         <= `TILE252.piton_pc_vld;
                  spc252_phy_pc_w          <= `TILE252.piton_pc;
                end
            end
    

            assign spc253_thread_id = 2'b00;
            assign spc253_rtl_pc = spc253_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(253*4)]   <= 1'b0;
                  active_thread[(253*4)+1] <= 1'b0;
                  active_thread[(253*4)+2] <= 1'b0;
                  active_thread[(253*4)+3] <= 1'b0;
                  spc253_inst_done         <= 0;
                  spc253_phy_pc_w          <= 0;
                end else begin
                  active_thread[(253*4)]   <= 1'b1;
                  active_thread[(253*4)+1] <= 1'b1;
                  active_thread[(253*4)+2] <= 1'b1;
                  active_thread[(253*4)+3] <= 1'b1;
                  spc253_inst_done         <= `TILE253.piton_pc_vld;
                  spc253_phy_pc_w          <= `TILE253.piton_pc;
                end
            end
    

            assign spc254_thread_id = 2'b00;
            assign spc254_rtl_pc = spc254_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(254*4)]   <= 1'b0;
                  active_thread[(254*4)+1] <= 1'b0;
                  active_thread[(254*4)+2] <= 1'b0;
                  active_thread[(254*4)+3] <= 1'b0;
                  spc254_inst_done         <= 0;
                  spc254_phy_pc_w          <= 0;
                end else begin
                  active_thread[(254*4)]   <= 1'b1;
                  active_thread[(254*4)+1] <= 1'b1;
                  active_thread[(254*4)+2] <= 1'b1;
                  active_thread[(254*4)+3] <= 1'b1;
                  spc254_inst_done         <= `TILE254.piton_pc_vld;
                  spc254_phy_pc_w          <= `TILE254.piton_pc;
                end
            end
    

            assign spc255_thread_id = 2'b00;
            assign spc255_rtl_pc = spc255_phy_pc_w;

            always @(posedge clk) begin
                if (~rst_l) begin
                  active_thread[(255*4)]   <= 1'b0;
                  active_thread[(255*4)+1] <= 1'b0;
                  active_thread[(255*4)+2] <= 1'b0;
                  active_thread[(255*4)+3] <= 1'b0;
                  spc255_inst_done         <= 0;
                  spc255_phy_pc_w          <= 0;
                end else begin
                  active_thread[(255*4)]   <= 1'b1;
                  active_thread[(255*4)+1] <= 1'b1;
                  active_thread[(255*4)+2] <= 1'b1;
                  active_thread[(255*4)+3] <= 1'b1;
                  spc255_inst_done         <= `TILE255.piton_pc_vld;
                  spc255_phy_pc_w          <= `TILE255.piton_pc;
                end
            end
    




reg           dummy;

task trap_extract;
    reg [2048:0] pc_str;
    reg [63:0]  tmp_val;
    integer     i;
    begin
        bad_trap_count = 0;

            if($value$plusargs("good_trap0=%h", tmp_val)) begin
                good_trap[0] = tmp_val;
                good_trap_exists[0] = 1'b1;
                //$display ("%t: good_trap %h", $time, good_trap[0]);
            end



            if($value$plusargs("bad_trap0=%h", tmp_val)) begin
                bad_trap[0] = tmp_val;
                bad_trap_exists[0] = 1'b1;
                //$display ("%t: bad_trap %h", $time, bad_trap[0]);
            end

        trap_count = good_trap_count > bad_trap_count ? good_trap_count :  bad_trap_count;

    end
endtask // trap_extract
// deceide pass or fail
integer       ind;
//post-silicon request
reg [63:0]    last_hit [31:0];
//indicate the 2nd time hit.
reg [31:0]    hitted;
initial hitted = 0;

reg first_rst;
initial begin
    //#20//need to wait for socket initializing.
     trap_extract;
    done    = 0;
    first_rst = 1;
    for(ind = 0;ind < `PITON_NUM_TILES; ind = ind + 1)timeout[ind] = 0;
end // initial begin
always @(posedge rst_l)begin
    if(first_rst)begin
        active_thread = 0;
        first_rst     = 0;
        done          = 0;
    end
end

task set_diag_done;
    input local_diag_done;

    begin
        if (local_diag_done) begin
            `TOP_MOD.diag_done = 1;
        end
    end
endtask


    wire[31:0] long_cpuid0;
    assign long_cpuid0 = {30'd0, spc0_thread_id};

    wire[31:0] long_cpuid1;
    assign long_cpuid1 = {30'd1, spc1_thread_id};

    wire[31:0] long_cpuid2;
    assign long_cpuid2 = {30'd2, spc2_thread_id};

    wire[31:0] long_cpuid3;
    assign long_cpuid3 = {30'd3, spc3_thread_id};

    wire[31:0] long_cpuid4;
    assign long_cpuid4 = {30'd4, spc4_thread_id};

    wire[31:0] long_cpuid5;
    assign long_cpuid5 = {30'd5, spc5_thread_id};

    wire[31:0] long_cpuid6;
    assign long_cpuid6 = {30'd6, spc6_thread_id};

    wire[31:0] long_cpuid7;
    assign long_cpuid7 = {30'd7, spc7_thread_id};

    wire[31:0] long_cpuid8;
    assign long_cpuid8 = {30'd8, spc8_thread_id};

    wire[31:0] long_cpuid9;
    assign long_cpuid9 = {30'd9, spc9_thread_id};

    wire[31:0] long_cpuid10;
    assign long_cpuid10 = {30'd10, spc10_thread_id};

    wire[31:0] long_cpuid11;
    assign long_cpuid11 = {30'd11, spc11_thread_id};

    wire[31:0] long_cpuid12;
    assign long_cpuid12 = {30'd12, spc12_thread_id};

    wire[31:0] long_cpuid13;
    assign long_cpuid13 = {30'd13, spc13_thread_id};

    wire[31:0] long_cpuid14;
    assign long_cpuid14 = {30'd14, spc14_thread_id};

    wire[31:0] long_cpuid15;
    assign long_cpuid15 = {30'd15, spc15_thread_id};

    wire[31:0] long_cpuid16;
    assign long_cpuid16 = {30'd16, spc16_thread_id};

    wire[31:0] long_cpuid17;
    assign long_cpuid17 = {30'd17, spc17_thread_id};

    wire[31:0] long_cpuid18;
    assign long_cpuid18 = {30'd18, spc18_thread_id};

    wire[31:0] long_cpuid19;
    assign long_cpuid19 = {30'd19, spc19_thread_id};

    wire[31:0] long_cpuid20;
    assign long_cpuid20 = {30'd20, spc20_thread_id};

    wire[31:0] long_cpuid21;
    assign long_cpuid21 = {30'd21, spc21_thread_id};

    wire[31:0] long_cpuid22;
    assign long_cpuid22 = {30'd22, spc22_thread_id};

    wire[31:0] long_cpuid23;
    assign long_cpuid23 = {30'd23, spc23_thread_id};

    wire[31:0] long_cpuid24;
    assign long_cpuid24 = {30'd24, spc24_thread_id};

    wire[31:0] long_cpuid25;
    assign long_cpuid25 = {30'd25, spc25_thread_id};

    wire[31:0] long_cpuid26;
    assign long_cpuid26 = {30'd26, spc26_thread_id};

    wire[31:0] long_cpuid27;
    assign long_cpuid27 = {30'd27, spc27_thread_id};

    wire[31:0] long_cpuid28;
    assign long_cpuid28 = {30'd28, spc28_thread_id};

    wire[31:0] long_cpuid29;
    assign long_cpuid29 = {30'd29, spc29_thread_id};

    wire[31:0] long_cpuid30;
    assign long_cpuid30 = {30'd30, spc30_thread_id};

    wire[31:0] long_cpuid31;
    assign long_cpuid31 = {30'd31, spc31_thread_id};

    wire[31:0] long_cpuid32;
    assign long_cpuid32 = {30'd32, spc32_thread_id};

    wire[31:0] long_cpuid33;
    assign long_cpuid33 = {30'd33, spc33_thread_id};

    wire[31:0] long_cpuid34;
    assign long_cpuid34 = {30'd34, spc34_thread_id};

    wire[31:0] long_cpuid35;
    assign long_cpuid35 = {30'd35, spc35_thread_id};

    wire[31:0] long_cpuid36;
    assign long_cpuid36 = {30'd36, spc36_thread_id};

    wire[31:0] long_cpuid37;
    assign long_cpuid37 = {30'd37, spc37_thread_id};

    wire[31:0] long_cpuid38;
    assign long_cpuid38 = {30'd38, spc38_thread_id};

    wire[31:0] long_cpuid39;
    assign long_cpuid39 = {30'd39, spc39_thread_id};

    wire[31:0] long_cpuid40;
    assign long_cpuid40 = {30'd40, spc40_thread_id};

    wire[31:0] long_cpuid41;
    assign long_cpuid41 = {30'd41, spc41_thread_id};

    wire[31:0] long_cpuid42;
    assign long_cpuid42 = {30'd42, spc42_thread_id};

    wire[31:0] long_cpuid43;
    assign long_cpuid43 = {30'd43, spc43_thread_id};

    wire[31:0] long_cpuid44;
    assign long_cpuid44 = {30'd44, spc44_thread_id};

    wire[31:0] long_cpuid45;
    assign long_cpuid45 = {30'd45, spc45_thread_id};

    wire[31:0] long_cpuid46;
    assign long_cpuid46 = {30'd46, spc46_thread_id};

    wire[31:0] long_cpuid47;
    assign long_cpuid47 = {30'd47, spc47_thread_id};

    wire[31:0] long_cpuid48;
    assign long_cpuid48 = {30'd48, spc48_thread_id};

    wire[31:0] long_cpuid49;
    assign long_cpuid49 = {30'd49, spc49_thread_id};

    wire[31:0] long_cpuid50;
    assign long_cpuid50 = {30'd50, spc50_thread_id};

    wire[31:0] long_cpuid51;
    assign long_cpuid51 = {30'd51, spc51_thread_id};

    wire[31:0] long_cpuid52;
    assign long_cpuid52 = {30'd52, spc52_thread_id};

    wire[31:0] long_cpuid53;
    assign long_cpuid53 = {30'd53, spc53_thread_id};

    wire[31:0] long_cpuid54;
    assign long_cpuid54 = {30'd54, spc54_thread_id};

    wire[31:0] long_cpuid55;
    assign long_cpuid55 = {30'd55, spc55_thread_id};

    wire[31:0] long_cpuid56;
    assign long_cpuid56 = {30'd56, spc56_thread_id};

    wire[31:0] long_cpuid57;
    assign long_cpuid57 = {30'd57, spc57_thread_id};

    wire[31:0] long_cpuid58;
    assign long_cpuid58 = {30'd58, spc58_thread_id};

    wire[31:0] long_cpuid59;
    assign long_cpuid59 = {30'd59, spc59_thread_id};

    wire[31:0] long_cpuid60;
    assign long_cpuid60 = {30'd60, spc60_thread_id};

    wire[31:0] long_cpuid61;
    assign long_cpuid61 = {30'd61, spc61_thread_id};

    wire[31:0] long_cpuid62;
    assign long_cpuid62 = {30'd62, spc62_thread_id};

    wire[31:0] long_cpuid63;
    assign long_cpuid63 = {30'd63, spc63_thread_id};

    wire[31:0] long_cpuid64;
    assign long_cpuid64 = {30'd64, spc64_thread_id};

    wire[31:0] long_cpuid65;
    assign long_cpuid65 = {30'd65, spc65_thread_id};

    wire[31:0] long_cpuid66;
    assign long_cpuid66 = {30'd66, spc66_thread_id};

    wire[31:0] long_cpuid67;
    assign long_cpuid67 = {30'd67, spc67_thread_id};

    wire[31:0] long_cpuid68;
    assign long_cpuid68 = {30'd68, spc68_thread_id};

    wire[31:0] long_cpuid69;
    assign long_cpuid69 = {30'd69, spc69_thread_id};

    wire[31:0] long_cpuid70;
    assign long_cpuid70 = {30'd70, spc70_thread_id};

    wire[31:0] long_cpuid71;
    assign long_cpuid71 = {30'd71, spc71_thread_id};

    wire[31:0] long_cpuid72;
    assign long_cpuid72 = {30'd72, spc72_thread_id};

    wire[31:0] long_cpuid73;
    assign long_cpuid73 = {30'd73, spc73_thread_id};

    wire[31:0] long_cpuid74;
    assign long_cpuid74 = {30'd74, spc74_thread_id};

    wire[31:0] long_cpuid75;
    assign long_cpuid75 = {30'd75, spc75_thread_id};

    wire[31:0] long_cpuid76;
    assign long_cpuid76 = {30'd76, spc76_thread_id};

    wire[31:0] long_cpuid77;
    assign long_cpuid77 = {30'd77, spc77_thread_id};

    wire[31:0] long_cpuid78;
    assign long_cpuid78 = {30'd78, spc78_thread_id};

    wire[31:0] long_cpuid79;
    assign long_cpuid79 = {30'd79, spc79_thread_id};

    wire[31:0] long_cpuid80;
    assign long_cpuid80 = {30'd80, spc80_thread_id};

    wire[31:0] long_cpuid81;
    assign long_cpuid81 = {30'd81, spc81_thread_id};

    wire[31:0] long_cpuid82;
    assign long_cpuid82 = {30'd82, spc82_thread_id};

    wire[31:0] long_cpuid83;
    assign long_cpuid83 = {30'd83, spc83_thread_id};

    wire[31:0] long_cpuid84;
    assign long_cpuid84 = {30'd84, spc84_thread_id};

    wire[31:0] long_cpuid85;
    assign long_cpuid85 = {30'd85, spc85_thread_id};

    wire[31:0] long_cpuid86;
    assign long_cpuid86 = {30'd86, spc86_thread_id};

    wire[31:0] long_cpuid87;
    assign long_cpuid87 = {30'd87, spc87_thread_id};

    wire[31:0] long_cpuid88;
    assign long_cpuid88 = {30'd88, spc88_thread_id};

    wire[31:0] long_cpuid89;
    assign long_cpuid89 = {30'd89, spc89_thread_id};

    wire[31:0] long_cpuid90;
    assign long_cpuid90 = {30'd90, spc90_thread_id};

    wire[31:0] long_cpuid91;
    assign long_cpuid91 = {30'd91, spc91_thread_id};

    wire[31:0] long_cpuid92;
    assign long_cpuid92 = {30'd92, spc92_thread_id};

    wire[31:0] long_cpuid93;
    assign long_cpuid93 = {30'd93, spc93_thread_id};

    wire[31:0] long_cpuid94;
    assign long_cpuid94 = {30'd94, spc94_thread_id};

    wire[31:0] long_cpuid95;
    assign long_cpuid95 = {30'd95, spc95_thread_id};

    wire[31:0] long_cpuid96;
    assign long_cpuid96 = {30'd96, spc96_thread_id};

    wire[31:0] long_cpuid97;
    assign long_cpuid97 = {30'd97, spc97_thread_id};

    wire[31:0] long_cpuid98;
    assign long_cpuid98 = {30'd98, spc98_thread_id};

    wire[31:0] long_cpuid99;
    assign long_cpuid99 = {30'd99, spc99_thread_id};

    wire[31:0] long_cpuid100;
    assign long_cpuid100 = {30'd100, spc100_thread_id};

    wire[31:0] long_cpuid101;
    assign long_cpuid101 = {30'd101, spc101_thread_id};

    wire[31:0] long_cpuid102;
    assign long_cpuid102 = {30'd102, spc102_thread_id};

    wire[31:0] long_cpuid103;
    assign long_cpuid103 = {30'd103, spc103_thread_id};

    wire[31:0] long_cpuid104;
    assign long_cpuid104 = {30'd104, spc104_thread_id};

    wire[31:0] long_cpuid105;
    assign long_cpuid105 = {30'd105, spc105_thread_id};

    wire[31:0] long_cpuid106;
    assign long_cpuid106 = {30'd106, spc106_thread_id};

    wire[31:0] long_cpuid107;
    assign long_cpuid107 = {30'd107, spc107_thread_id};

    wire[31:0] long_cpuid108;
    assign long_cpuid108 = {30'd108, spc108_thread_id};

    wire[31:0] long_cpuid109;
    assign long_cpuid109 = {30'd109, spc109_thread_id};

    wire[31:0] long_cpuid110;
    assign long_cpuid110 = {30'd110, spc110_thread_id};

    wire[31:0] long_cpuid111;
    assign long_cpuid111 = {30'd111, spc111_thread_id};

    wire[31:0] long_cpuid112;
    assign long_cpuid112 = {30'd112, spc112_thread_id};

    wire[31:0] long_cpuid113;
    assign long_cpuid113 = {30'd113, spc113_thread_id};

    wire[31:0] long_cpuid114;
    assign long_cpuid114 = {30'd114, spc114_thread_id};

    wire[31:0] long_cpuid115;
    assign long_cpuid115 = {30'd115, spc115_thread_id};

    wire[31:0] long_cpuid116;
    assign long_cpuid116 = {30'd116, spc116_thread_id};

    wire[31:0] long_cpuid117;
    assign long_cpuid117 = {30'd117, spc117_thread_id};

    wire[31:0] long_cpuid118;
    assign long_cpuid118 = {30'd118, spc118_thread_id};

    wire[31:0] long_cpuid119;
    assign long_cpuid119 = {30'd119, spc119_thread_id};

    wire[31:0] long_cpuid120;
    assign long_cpuid120 = {30'd120, spc120_thread_id};

    wire[31:0] long_cpuid121;
    assign long_cpuid121 = {30'd121, spc121_thread_id};

    wire[31:0] long_cpuid122;
    assign long_cpuid122 = {30'd122, spc122_thread_id};

    wire[31:0] long_cpuid123;
    assign long_cpuid123 = {30'd123, spc123_thread_id};

    wire[31:0] long_cpuid124;
    assign long_cpuid124 = {30'd124, spc124_thread_id};

    wire[31:0] long_cpuid125;
    assign long_cpuid125 = {30'd125, spc125_thread_id};

    wire[31:0] long_cpuid126;
    assign long_cpuid126 = {30'd126, spc126_thread_id};

    wire[31:0] long_cpuid127;
    assign long_cpuid127 = {30'd127, spc127_thread_id};

    wire[31:0] long_cpuid128;
    assign long_cpuid128 = {30'd128, spc128_thread_id};

    wire[31:0] long_cpuid129;
    assign long_cpuid129 = {30'd129, spc129_thread_id};

    wire[31:0] long_cpuid130;
    assign long_cpuid130 = {30'd130, spc130_thread_id};

    wire[31:0] long_cpuid131;
    assign long_cpuid131 = {30'd131, spc131_thread_id};

    wire[31:0] long_cpuid132;
    assign long_cpuid132 = {30'd132, spc132_thread_id};

    wire[31:0] long_cpuid133;
    assign long_cpuid133 = {30'd133, spc133_thread_id};

    wire[31:0] long_cpuid134;
    assign long_cpuid134 = {30'd134, spc134_thread_id};

    wire[31:0] long_cpuid135;
    assign long_cpuid135 = {30'd135, spc135_thread_id};

    wire[31:0] long_cpuid136;
    assign long_cpuid136 = {30'd136, spc136_thread_id};

    wire[31:0] long_cpuid137;
    assign long_cpuid137 = {30'd137, spc137_thread_id};

    wire[31:0] long_cpuid138;
    assign long_cpuid138 = {30'd138, spc138_thread_id};

    wire[31:0] long_cpuid139;
    assign long_cpuid139 = {30'd139, spc139_thread_id};

    wire[31:0] long_cpuid140;
    assign long_cpuid140 = {30'd140, spc140_thread_id};

    wire[31:0] long_cpuid141;
    assign long_cpuid141 = {30'd141, spc141_thread_id};

    wire[31:0] long_cpuid142;
    assign long_cpuid142 = {30'd142, spc142_thread_id};

    wire[31:0] long_cpuid143;
    assign long_cpuid143 = {30'd143, spc143_thread_id};

    wire[31:0] long_cpuid144;
    assign long_cpuid144 = {30'd144, spc144_thread_id};

    wire[31:0] long_cpuid145;
    assign long_cpuid145 = {30'd145, spc145_thread_id};

    wire[31:0] long_cpuid146;
    assign long_cpuid146 = {30'd146, spc146_thread_id};

    wire[31:0] long_cpuid147;
    assign long_cpuid147 = {30'd147, spc147_thread_id};

    wire[31:0] long_cpuid148;
    assign long_cpuid148 = {30'd148, spc148_thread_id};

    wire[31:0] long_cpuid149;
    assign long_cpuid149 = {30'd149, spc149_thread_id};

    wire[31:0] long_cpuid150;
    assign long_cpuid150 = {30'd150, spc150_thread_id};

    wire[31:0] long_cpuid151;
    assign long_cpuid151 = {30'd151, spc151_thread_id};

    wire[31:0] long_cpuid152;
    assign long_cpuid152 = {30'd152, spc152_thread_id};

    wire[31:0] long_cpuid153;
    assign long_cpuid153 = {30'd153, spc153_thread_id};

    wire[31:0] long_cpuid154;
    assign long_cpuid154 = {30'd154, spc154_thread_id};

    wire[31:0] long_cpuid155;
    assign long_cpuid155 = {30'd155, spc155_thread_id};

    wire[31:0] long_cpuid156;
    assign long_cpuid156 = {30'd156, spc156_thread_id};

    wire[31:0] long_cpuid157;
    assign long_cpuid157 = {30'd157, spc157_thread_id};

    wire[31:0] long_cpuid158;
    assign long_cpuid158 = {30'd158, spc158_thread_id};

    wire[31:0] long_cpuid159;
    assign long_cpuid159 = {30'd159, spc159_thread_id};

    wire[31:0] long_cpuid160;
    assign long_cpuid160 = {30'd160, spc160_thread_id};

    wire[31:0] long_cpuid161;
    assign long_cpuid161 = {30'd161, spc161_thread_id};

    wire[31:0] long_cpuid162;
    assign long_cpuid162 = {30'd162, spc162_thread_id};

    wire[31:0] long_cpuid163;
    assign long_cpuid163 = {30'd163, spc163_thread_id};

    wire[31:0] long_cpuid164;
    assign long_cpuid164 = {30'd164, spc164_thread_id};

    wire[31:0] long_cpuid165;
    assign long_cpuid165 = {30'd165, spc165_thread_id};

    wire[31:0] long_cpuid166;
    assign long_cpuid166 = {30'd166, spc166_thread_id};

    wire[31:0] long_cpuid167;
    assign long_cpuid167 = {30'd167, spc167_thread_id};

    wire[31:0] long_cpuid168;
    assign long_cpuid168 = {30'd168, spc168_thread_id};

    wire[31:0] long_cpuid169;
    assign long_cpuid169 = {30'd169, spc169_thread_id};

    wire[31:0] long_cpuid170;
    assign long_cpuid170 = {30'd170, spc170_thread_id};

    wire[31:0] long_cpuid171;
    assign long_cpuid171 = {30'd171, spc171_thread_id};

    wire[31:0] long_cpuid172;
    assign long_cpuid172 = {30'd172, spc172_thread_id};

    wire[31:0] long_cpuid173;
    assign long_cpuid173 = {30'd173, spc173_thread_id};

    wire[31:0] long_cpuid174;
    assign long_cpuid174 = {30'd174, spc174_thread_id};

    wire[31:0] long_cpuid175;
    assign long_cpuid175 = {30'd175, spc175_thread_id};

    wire[31:0] long_cpuid176;
    assign long_cpuid176 = {30'd176, spc176_thread_id};

    wire[31:0] long_cpuid177;
    assign long_cpuid177 = {30'd177, spc177_thread_id};

    wire[31:0] long_cpuid178;
    assign long_cpuid178 = {30'd178, spc178_thread_id};

    wire[31:0] long_cpuid179;
    assign long_cpuid179 = {30'd179, spc179_thread_id};

    wire[31:0] long_cpuid180;
    assign long_cpuid180 = {30'd180, spc180_thread_id};

    wire[31:0] long_cpuid181;
    assign long_cpuid181 = {30'd181, spc181_thread_id};

    wire[31:0] long_cpuid182;
    assign long_cpuid182 = {30'd182, spc182_thread_id};

    wire[31:0] long_cpuid183;
    assign long_cpuid183 = {30'd183, spc183_thread_id};

    wire[31:0] long_cpuid184;
    assign long_cpuid184 = {30'd184, spc184_thread_id};

    wire[31:0] long_cpuid185;
    assign long_cpuid185 = {30'd185, spc185_thread_id};

    wire[31:0] long_cpuid186;
    assign long_cpuid186 = {30'd186, spc186_thread_id};

    wire[31:0] long_cpuid187;
    assign long_cpuid187 = {30'd187, spc187_thread_id};

    wire[31:0] long_cpuid188;
    assign long_cpuid188 = {30'd188, spc188_thread_id};

    wire[31:0] long_cpuid189;
    assign long_cpuid189 = {30'd189, spc189_thread_id};

    wire[31:0] long_cpuid190;
    assign long_cpuid190 = {30'd190, spc190_thread_id};

    wire[31:0] long_cpuid191;
    assign long_cpuid191 = {30'd191, spc191_thread_id};

    wire[31:0] long_cpuid192;
    assign long_cpuid192 = {30'd192, spc192_thread_id};

    wire[31:0] long_cpuid193;
    assign long_cpuid193 = {30'd193, spc193_thread_id};

    wire[31:0] long_cpuid194;
    assign long_cpuid194 = {30'd194, spc194_thread_id};

    wire[31:0] long_cpuid195;
    assign long_cpuid195 = {30'd195, spc195_thread_id};

    wire[31:0] long_cpuid196;
    assign long_cpuid196 = {30'd196, spc196_thread_id};

    wire[31:0] long_cpuid197;
    assign long_cpuid197 = {30'd197, spc197_thread_id};

    wire[31:0] long_cpuid198;
    assign long_cpuid198 = {30'd198, spc198_thread_id};

    wire[31:0] long_cpuid199;
    assign long_cpuid199 = {30'd199, spc199_thread_id};

    wire[31:0] long_cpuid200;
    assign long_cpuid200 = {30'd200, spc200_thread_id};

    wire[31:0] long_cpuid201;
    assign long_cpuid201 = {30'd201, spc201_thread_id};

    wire[31:0] long_cpuid202;
    assign long_cpuid202 = {30'd202, spc202_thread_id};

    wire[31:0] long_cpuid203;
    assign long_cpuid203 = {30'd203, spc203_thread_id};

    wire[31:0] long_cpuid204;
    assign long_cpuid204 = {30'd204, spc204_thread_id};

    wire[31:0] long_cpuid205;
    assign long_cpuid205 = {30'd205, spc205_thread_id};

    wire[31:0] long_cpuid206;
    assign long_cpuid206 = {30'd206, spc206_thread_id};

    wire[31:0] long_cpuid207;
    assign long_cpuid207 = {30'd207, spc207_thread_id};

    wire[31:0] long_cpuid208;
    assign long_cpuid208 = {30'd208, spc208_thread_id};

    wire[31:0] long_cpuid209;
    assign long_cpuid209 = {30'd209, spc209_thread_id};

    wire[31:0] long_cpuid210;
    assign long_cpuid210 = {30'd210, spc210_thread_id};

    wire[31:0] long_cpuid211;
    assign long_cpuid211 = {30'd211, spc211_thread_id};

    wire[31:0] long_cpuid212;
    assign long_cpuid212 = {30'd212, spc212_thread_id};

    wire[31:0] long_cpuid213;
    assign long_cpuid213 = {30'd213, spc213_thread_id};

    wire[31:0] long_cpuid214;
    assign long_cpuid214 = {30'd214, spc214_thread_id};

    wire[31:0] long_cpuid215;
    assign long_cpuid215 = {30'd215, spc215_thread_id};

    wire[31:0] long_cpuid216;
    assign long_cpuid216 = {30'd216, spc216_thread_id};

    wire[31:0] long_cpuid217;
    assign long_cpuid217 = {30'd217, spc217_thread_id};

    wire[31:0] long_cpuid218;
    assign long_cpuid218 = {30'd218, spc218_thread_id};

    wire[31:0] long_cpuid219;
    assign long_cpuid219 = {30'd219, spc219_thread_id};

    wire[31:0] long_cpuid220;
    assign long_cpuid220 = {30'd220, spc220_thread_id};

    wire[31:0] long_cpuid221;
    assign long_cpuid221 = {30'd221, spc221_thread_id};

    wire[31:0] long_cpuid222;
    assign long_cpuid222 = {30'd222, spc222_thread_id};

    wire[31:0] long_cpuid223;
    assign long_cpuid223 = {30'd223, spc223_thread_id};

    wire[31:0] long_cpuid224;
    assign long_cpuid224 = {30'd224, spc224_thread_id};

    wire[31:0] long_cpuid225;
    assign long_cpuid225 = {30'd225, spc225_thread_id};

    wire[31:0] long_cpuid226;
    assign long_cpuid226 = {30'd226, spc226_thread_id};

    wire[31:0] long_cpuid227;
    assign long_cpuid227 = {30'd227, spc227_thread_id};

    wire[31:0] long_cpuid228;
    assign long_cpuid228 = {30'd228, spc228_thread_id};

    wire[31:0] long_cpuid229;
    assign long_cpuid229 = {30'd229, spc229_thread_id};

    wire[31:0] long_cpuid230;
    assign long_cpuid230 = {30'd230, spc230_thread_id};

    wire[31:0] long_cpuid231;
    assign long_cpuid231 = {30'd231, spc231_thread_id};

    wire[31:0] long_cpuid232;
    assign long_cpuid232 = {30'd232, spc232_thread_id};

    wire[31:0] long_cpuid233;
    assign long_cpuid233 = {30'd233, spc233_thread_id};

    wire[31:0] long_cpuid234;
    assign long_cpuid234 = {30'd234, spc234_thread_id};

    wire[31:0] long_cpuid235;
    assign long_cpuid235 = {30'd235, spc235_thread_id};

    wire[31:0] long_cpuid236;
    assign long_cpuid236 = {30'd236, spc236_thread_id};

    wire[31:0] long_cpuid237;
    assign long_cpuid237 = {30'd237, spc237_thread_id};

    wire[31:0] long_cpuid238;
    assign long_cpuid238 = {30'd238, spc238_thread_id};

    wire[31:0] long_cpuid239;
    assign long_cpuid239 = {30'd239, spc239_thread_id};

    wire[31:0] long_cpuid240;
    assign long_cpuid240 = {30'd240, spc240_thread_id};

    wire[31:0] long_cpuid241;
    assign long_cpuid241 = {30'd241, spc241_thread_id};

    wire[31:0] long_cpuid242;
    assign long_cpuid242 = {30'd242, spc242_thread_id};

    wire[31:0] long_cpuid243;
    assign long_cpuid243 = {30'd243, spc243_thread_id};

    wire[31:0] long_cpuid244;
    assign long_cpuid244 = {30'd244, spc244_thread_id};

    wire[31:0] long_cpuid245;
    assign long_cpuid245 = {30'd245, spc245_thread_id};

    wire[31:0] long_cpuid246;
    assign long_cpuid246 = {30'd246, spc246_thread_id};

    wire[31:0] long_cpuid247;
    assign long_cpuid247 = {30'd247, spc247_thread_id};

    wire[31:0] long_cpuid248;
    assign long_cpuid248 = {30'd248, spc248_thread_id};

    wire[31:0] long_cpuid249;
    assign long_cpuid249 = {30'd249, spc249_thread_id};

    wire[31:0] long_cpuid250;
    assign long_cpuid250 = {30'd250, spc250_thread_id};

    wire[31:0] long_cpuid251;
    assign long_cpuid251 = {30'd251, spc251_thread_id};

    wire[31:0] long_cpuid252;
    assign long_cpuid252 = {30'd252, spc252_thread_id};

    wire[31:0] long_cpuid253;
    assign long_cpuid253 = {30'd253, spc253_thread_id};

    wire[31:0] long_cpuid254;
    assign long_cpuid254 = {30'd254, spc254_thread_id};

    wire[31:0] long_cpuid255;
    assign long_cpuid255 = {30'd255, spc255_thread_id};


always @* begin
done[0]   = spc0_inst_done;//sparc 0
done[1]   = spc1_inst_done;//sparc 1
done[2]   = spc2_inst_done;//sparc 2
done[3]   = spc3_inst_done;//sparc 3
done[4]   = spc4_inst_done;//sparc 4
done[5]   = spc5_inst_done;//sparc 5
done[6]   = spc6_inst_done;//sparc 6
done[7]   = spc7_inst_done;//sparc 7
done[8]   = spc8_inst_done;//sparc 8
done[9]   = spc9_inst_done;//sparc 9
done[10]   = spc10_inst_done;//sparc 10
done[11]   = spc11_inst_done;//sparc 11
done[12]   = spc12_inst_done;//sparc 12
done[13]   = spc13_inst_done;//sparc 13
done[14]   = spc14_inst_done;//sparc 14
done[15]   = spc15_inst_done;//sparc 15
done[16]   = spc16_inst_done;//sparc 16
done[17]   = spc17_inst_done;//sparc 17
done[18]   = spc18_inst_done;//sparc 18
done[19]   = spc19_inst_done;//sparc 19
done[20]   = spc20_inst_done;//sparc 20
done[21]   = spc21_inst_done;//sparc 21
done[22]   = spc22_inst_done;//sparc 22
done[23]   = spc23_inst_done;//sparc 23
done[24]   = spc24_inst_done;//sparc 24
done[25]   = spc25_inst_done;//sparc 25
done[26]   = spc26_inst_done;//sparc 26
done[27]   = spc27_inst_done;//sparc 27
done[28]   = spc28_inst_done;//sparc 28
done[29]   = spc29_inst_done;//sparc 29
done[30]   = spc30_inst_done;//sparc 30
done[31]   = spc31_inst_done;//sparc 31
done[32]   = spc32_inst_done;//sparc 32
done[33]   = spc33_inst_done;//sparc 33
done[34]   = spc34_inst_done;//sparc 34
done[35]   = spc35_inst_done;//sparc 35
done[36]   = spc36_inst_done;//sparc 36
done[37]   = spc37_inst_done;//sparc 37
done[38]   = spc38_inst_done;//sparc 38
done[39]   = spc39_inst_done;//sparc 39
done[40]   = spc40_inst_done;//sparc 40
done[41]   = spc41_inst_done;//sparc 41
done[42]   = spc42_inst_done;//sparc 42
done[43]   = spc43_inst_done;//sparc 43
done[44]   = spc44_inst_done;//sparc 44
done[45]   = spc45_inst_done;//sparc 45
done[46]   = spc46_inst_done;//sparc 46
done[47]   = spc47_inst_done;//sparc 47
done[48]   = spc48_inst_done;//sparc 48
done[49]   = spc49_inst_done;//sparc 49
done[50]   = spc50_inst_done;//sparc 50
done[51]   = spc51_inst_done;//sparc 51
done[52]   = spc52_inst_done;//sparc 52
done[53]   = spc53_inst_done;//sparc 53
done[54]   = spc54_inst_done;//sparc 54
done[55]   = spc55_inst_done;//sparc 55
done[56]   = spc56_inst_done;//sparc 56
done[57]   = spc57_inst_done;//sparc 57
done[58]   = spc58_inst_done;//sparc 58
done[59]   = spc59_inst_done;//sparc 59
done[60]   = spc60_inst_done;//sparc 60
done[61]   = spc61_inst_done;//sparc 61
done[62]   = spc62_inst_done;//sparc 62
done[63]   = spc63_inst_done;//sparc 63
done[64]   = spc64_inst_done;//sparc 64
done[65]   = spc65_inst_done;//sparc 65
done[66]   = spc66_inst_done;//sparc 66
done[67]   = spc67_inst_done;//sparc 67
done[68]   = spc68_inst_done;//sparc 68
done[69]   = spc69_inst_done;//sparc 69
done[70]   = spc70_inst_done;//sparc 70
done[71]   = spc71_inst_done;//sparc 71
done[72]   = spc72_inst_done;//sparc 72
done[73]   = spc73_inst_done;//sparc 73
done[74]   = spc74_inst_done;//sparc 74
done[75]   = spc75_inst_done;//sparc 75
done[76]   = spc76_inst_done;//sparc 76
done[77]   = spc77_inst_done;//sparc 77
done[78]   = spc78_inst_done;//sparc 78
done[79]   = spc79_inst_done;//sparc 79
done[80]   = spc80_inst_done;//sparc 80
done[81]   = spc81_inst_done;//sparc 81
done[82]   = spc82_inst_done;//sparc 82
done[83]   = spc83_inst_done;//sparc 83
done[84]   = spc84_inst_done;//sparc 84
done[85]   = spc85_inst_done;//sparc 85
done[86]   = spc86_inst_done;//sparc 86
done[87]   = spc87_inst_done;//sparc 87
done[88]   = spc88_inst_done;//sparc 88
done[89]   = spc89_inst_done;//sparc 89
done[90]   = spc90_inst_done;//sparc 90
done[91]   = spc91_inst_done;//sparc 91
done[92]   = spc92_inst_done;//sparc 92
done[93]   = spc93_inst_done;//sparc 93
done[94]   = spc94_inst_done;//sparc 94
done[95]   = spc95_inst_done;//sparc 95
done[96]   = spc96_inst_done;//sparc 96
done[97]   = spc97_inst_done;//sparc 97
done[98]   = spc98_inst_done;//sparc 98
done[99]   = spc99_inst_done;//sparc 99
done[100]   = spc100_inst_done;//sparc 100
done[101]   = spc101_inst_done;//sparc 101
done[102]   = spc102_inst_done;//sparc 102
done[103]   = spc103_inst_done;//sparc 103
done[104]   = spc104_inst_done;//sparc 104
done[105]   = spc105_inst_done;//sparc 105
done[106]   = spc106_inst_done;//sparc 106
done[107]   = spc107_inst_done;//sparc 107
done[108]   = spc108_inst_done;//sparc 108
done[109]   = spc109_inst_done;//sparc 109
done[110]   = spc110_inst_done;//sparc 110
done[111]   = spc111_inst_done;//sparc 111
done[112]   = spc112_inst_done;//sparc 112
done[113]   = spc113_inst_done;//sparc 113
done[114]   = spc114_inst_done;//sparc 114
done[115]   = spc115_inst_done;//sparc 115
done[116]   = spc116_inst_done;//sparc 116
done[117]   = spc117_inst_done;//sparc 117
done[118]   = spc118_inst_done;//sparc 118
done[119]   = spc119_inst_done;//sparc 119
done[120]   = spc120_inst_done;//sparc 120
done[121]   = spc121_inst_done;//sparc 121
done[122]   = spc122_inst_done;//sparc 122
done[123]   = spc123_inst_done;//sparc 123
done[124]   = spc124_inst_done;//sparc 124
done[125]   = spc125_inst_done;//sparc 125
done[126]   = spc126_inst_done;//sparc 126
done[127]   = spc127_inst_done;//sparc 127
done[128]   = spc128_inst_done;//sparc 128
done[129]   = spc129_inst_done;//sparc 129
done[130]   = spc130_inst_done;//sparc 130
done[131]   = spc131_inst_done;//sparc 131
done[132]   = spc132_inst_done;//sparc 132
done[133]   = spc133_inst_done;//sparc 133
done[134]   = spc134_inst_done;//sparc 134
done[135]   = spc135_inst_done;//sparc 135
done[136]   = spc136_inst_done;//sparc 136
done[137]   = spc137_inst_done;//sparc 137
done[138]   = spc138_inst_done;//sparc 138
done[139]   = spc139_inst_done;//sparc 139
done[140]   = spc140_inst_done;//sparc 140
done[141]   = spc141_inst_done;//sparc 141
done[142]   = spc142_inst_done;//sparc 142
done[143]   = spc143_inst_done;//sparc 143
done[144]   = spc144_inst_done;//sparc 144
done[145]   = spc145_inst_done;//sparc 145
done[146]   = spc146_inst_done;//sparc 146
done[147]   = spc147_inst_done;//sparc 147
done[148]   = spc148_inst_done;//sparc 148
done[149]   = spc149_inst_done;//sparc 149
done[150]   = spc150_inst_done;//sparc 150
done[151]   = spc151_inst_done;//sparc 151
done[152]   = spc152_inst_done;//sparc 152
done[153]   = spc153_inst_done;//sparc 153
done[154]   = spc154_inst_done;//sparc 154
done[155]   = spc155_inst_done;//sparc 155
done[156]   = spc156_inst_done;//sparc 156
done[157]   = spc157_inst_done;//sparc 157
done[158]   = spc158_inst_done;//sparc 158
done[159]   = spc159_inst_done;//sparc 159
done[160]   = spc160_inst_done;//sparc 160
done[161]   = spc161_inst_done;//sparc 161
done[162]   = spc162_inst_done;//sparc 162
done[163]   = spc163_inst_done;//sparc 163
done[164]   = spc164_inst_done;//sparc 164
done[165]   = spc165_inst_done;//sparc 165
done[166]   = spc166_inst_done;//sparc 166
done[167]   = spc167_inst_done;//sparc 167
done[168]   = spc168_inst_done;//sparc 168
done[169]   = spc169_inst_done;//sparc 169
done[170]   = spc170_inst_done;//sparc 170
done[171]   = spc171_inst_done;//sparc 171
done[172]   = spc172_inst_done;//sparc 172
done[173]   = spc173_inst_done;//sparc 173
done[174]   = spc174_inst_done;//sparc 174
done[175]   = spc175_inst_done;//sparc 175
done[176]   = spc176_inst_done;//sparc 176
done[177]   = spc177_inst_done;//sparc 177
done[178]   = spc178_inst_done;//sparc 178
done[179]   = spc179_inst_done;//sparc 179
done[180]   = spc180_inst_done;//sparc 180
done[181]   = spc181_inst_done;//sparc 181
done[182]   = spc182_inst_done;//sparc 182
done[183]   = spc183_inst_done;//sparc 183
done[184]   = spc184_inst_done;//sparc 184
done[185]   = spc185_inst_done;//sparc 185
done[186]   = spc186_inst_done;//sparc 186
done[187]   = spc187_inst_done;//sparc 187
done[188]   = spc188_inst_done;//sparc 188
done[189]   = spc189_inst_done;//sparc 189
done[190]   = spc190_inst_done;//sparc 190
done[191]   = spc191_inst_done;//sparc 191
done[192]   = spc192_inst_done;//sparc 192
done[193]   = spc193_inst_done;//sparc 193
done[194]   = spc194_inst_done;//sparc 194
done[195]   = spc195_inst_done;//sparc 195
done[196]   = spc196_inst_done;//sparc 196
done[197]   = spc197_inst_done;//sparc 197
done[198]   = spc198_inst_done;//sparc 198
done[199]   = spc199_inst_done;//sparc 199
done[200]   = spc200_inst_done;//sparc 200
done[201]   = spc201_inst_done;//sparc 201
done[202]   = spc202_inst_done;//sparc 202
done[203]   = spc203_inst_done;//sparc 203
done[204]   = spc204_inst_done;//sparc 204
done[205]   = spc205_inst_done;//sparc 205
done[206]   = spc206_inst_done;//sparc 206
done[207]   = spc207_inst_done;//sparc 207
done[208]   = spc208_inst_done;//sparc 208
done[209]   = spc209_inst_done;//sparc 209
done[210]   = spc210_inst_done;//sparc 210
done[211]   = spc211_inst_done;//sparc 211
done[212]   = spc212_inst_done;//sparc 212
done[213]   = spc213_inst_done;//sparc 213
done[214]   = spc214_inst_done;//sparc 214
done[215]   = spc215_inst_done;//sparc 215
done[216]   = spc216_inst_done;//sparc 216
done[217]   = spc217_inst_done;//sparc 217
done[218]   = spc218_inst_done;//sparc 218
done[219]   = spc219_inst_done;//sparc 219
done[220]   = spc220_inst_done;//sparc 220
done[221]   = spc221_inst_done;//sparc 221
done[222]   = spc222_inst_done;//sparc 222
done[223]   = spc223_inst_done;//sparc 223
done[224]   = spc224_inst_done;//sparc 224
done[225]   = spc225_inst_done;//sparc 225
done[226]   = spc226_inst_done;//sparc 226
done[227]   = spc227_inst_done;//sparc 227
done[228]   = spc228_inst_done;//sparc 228
done[229]   = spc229_inst_done;//sparc 229
done[230]   = spc230_inst_done;//sparc 230
done[231]   = spc231_inst_done;//sparc 231
done[232]   = spc232_inst_done;//sparc 232
done[233]   = spc233_inst_done;//sparc 233
done[234]   = spc234_inst_done;//sparc 234
done[235]   = spc235_inst_done;//sparc 235
done[236]   = spc236_inst_done;//sparc 236
done[237]   = spc237_inst_done;//sparc 237
done[238]   = spc238_inst_done;//sparc 238
done[239]   = spc239_inst_done;//sparc 239
done[240]   = spc240_inst_done;//sparc 240
done[241]   = spc241_inst_done;//sparc 241
done[242]   = spc242_inst_done;//sparc 242
done[243]   = spc243_inst_done;//sparc 243
done[244]   = spc244_inst_done;//sparc 244
done[245]   = spc245_inst_done;//sparc 245
done[246]   = spc246_inst_done;//sparc 246
done[247]   = spc247_inst_done;//sparc 247
done[248]   = spc248_inst_done;//sparc 248
done[249]   = spc249_inst_done;//sparc 249
done[250]   = spc250_inst_done;//sparc 250
done[251]   = spc251_inst_done;//sparc 251
done[252]   = spc252_inst_done;//sparc 252
done[253]   = spc253_inst_done;//sparc 253
done[254]   = spc254_inst_done;//sparc 254
done[255]   = spc255_inst_done;//sparc 255


end



string linebuf0 = "";
logic hitMadPrint0 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc0_inst_done && ((spc0_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint0 = 1;
       linebuf0 = {linebuf0, spc0_phy_pc_w[8:1]};
       if (spc0_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 0, linebuf0);
          linebuf0 = "";
       end
    end else begin
       hitMadPrint0 = 0;
    end
  end
end


string linebuf1 = "";
logic hitMadPrint1 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc1_inst_done && ((spc1_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint1 = 1;
       linebuf1 = {linebuf1, spc1_phy_pc_w[8:1]};
       if (spc1_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 1, linebuf1);
          linebuf1 = "";
       end
    end else begin
       hitMadPrint1 = 0;
    end
  end
end


string linebuf2 = "";
logic hitMadPrint2 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc2_inst_done && ((spc2_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint2 = 1;
       linebuf2 = {linebuf2, spc2_phy_pc_w[8:1]};
       if (spc2_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 2, linebuf2);
          linebuf2 = "";
       end
    end else begin
       hitMadPrint2 = 0;
    end
  end
end


string linebuf3 = "";
logic hitMadPrint3 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc3_inst_done && ((spc3_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint3 = 1;
       linebuf3 = {linebuf3, spc3_phy_pc_w[8:1]};
       if (spc3_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 3, linebuf3);
          linebuf3 = "";
       end
    end else begin
       hitMadPrint3 = 0;
    end
  end
end


string linebuf4 = "";
logic hitMadPrint4 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc4_inst_done && ((spc4_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint4 = 1;
       linebuf4 = {linebuf4, spc4_phy_pc_w[8:1]};
       if (spc4_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 4, linebuf4);
          linebuf4 = "";
       end
    end else begin
       hitMadPrint4 = 0;
    end
  end
end


string linebuf5 = "";
logic hitMadPrint5 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc5_inst_done && ((spc5_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint5 = 1;
       linebuf5 = {linebuf5, spc5_phy_pc_w[8:1]};
       if (spc5_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 5, linebuf5);
          linebuf5 = "";
       end
    end else begin
       hitMadPrint5 = 0;
    end
  end
end


string linebuf6 = "";
logic hitMadPrint6 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc6_inst_done && ((spc6_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint6 = 1;
       linebuf6 = {linebuf6, spc6_phy_pc_w[8:1]};
       if (spc6_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 6, linebuf6);
          linebuf6 = "";
       end
    end else begin
       hitMadPrint6 = 0;
    end
  end
end


string linebuf7 = "";
logic hitMadPrint7 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc7_inst_done && ((spc7_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint7 = 1;
       linebuf7 = {linebuf7, spc7_phy_pc_w[8:1]};
       if (spc7_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 7, linebuf7);
          linebuf7 = "";
       end
    end else begin
       hitMadPrint7 = 0;
    end
  end
end


string linebuf8 = "";
logic hitMadPrint8 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc8_inst_done && ((spc8_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint8 = 1;
       linebuf8 = {linebuf8, spc8_phy_pc_w[8:1]};
       if (spc8_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 8, linebuf8);
          linebuf8 = "";
       end
    end else begin
       hitMadPrint8 = 0;
    end
  end
end


string linebuf9 = "";
logic hitMadPrint9 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc9_inst_done && ((spc9_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint9 = 1;
       linebuf9 = {linebuf9, spc9_phy_pc_w[8:1]};
       if (spc9_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 9, linebuf9);
          linebuf9 = "";
       end
    end else begin
       hitMadPrint9 = 0;
    end
  end
end


string linebuf10 = "";
logic hitMadPrint10 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc10_inst_done && ((spc10_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint10 = 1;
       linebuf10 = {linebuf10, spc10_phy_pc_w[8:1]};
       if (spc10_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 10, linebuf10);
          linebuf10 = "";
       end
    end else begin
       hitMadPrint10 = 0;
    end
  end
end


string linebuf11 = "";
logic hitMadPrint11 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc11_inst_done && ((spc11_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint11 = 1;
       linebuf11 = {linebuf11, spc11_phy_pc_w[8:1]};
       if (spc11_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 11, linebuf11);
          linebuf11 = "";
       end
    end else begin
       hitMadPrint11 = 0;
    end
  end
end


string linebuf12 = "";
logic hitMadPrint12 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc12_inst_done && ((spc12_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint12 = 1;
       linebuf12 = {linebuf12, spc12_phy_pc_w[8:1]};
       if (spc12_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 12, linebuf12);
          linebuf12 = "";
       end
    end else begin
       hitMadPrint12 = 0;
    end
  end
end


string linebuf13 = "";
logic hitMadPrint13 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc13_inst_done && ((spc13_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint13 = 1;
       linebuf13 = {linebuf13, spc13_phy_pc_w[8:1]};
       if (spc13_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 13, linebuf13);
          linebuf13 = "";
       end
    end else begin
       hitMadPrint13 = 0;
    end
  end
end


string linebuf14 = "";
logic hitMadPrint14 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc14_inst_done && ((spc14_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint14 = 1;
       linebuf14 = {linebuf14, spc14_phy_pc_w[8:1]};
       if (spc14_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 14, linebuf14);
          linebuf14 = "";
       end
    end else begin
       hitMadPrint14 = 0;
    end
  end
end


string linebuf15 = "";
logic hitMadPrint15 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc15_inst_done && ((spc15_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint15 = 1;
       linebuf15 = {linebuf15, spc15_phy_pc_w[8:1]};
       if (spc15_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 15, linebuf15);
          linebuf15 = "";
       end
    end else begin
       hitMadPrint15 = 0;
    end
  end
end


string linebuf16 = "";
logic hitMadPrint16 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc16_inst_done && ((spc16_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint16 = 1;
       linebuf16 = {linebuf16, spc16_phy_pc_w[8:1]};
       if (spc16_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 16, linebuf16);
          linebuf16 = "";
       end
    end else begin
       hitMadPrint16 = 0;
    end
  end
end


string linebuf17 = "";
logic hitMadPrint17 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc17_inst_done && ((spc17_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint17 = 1;
       linebuf17 = {linebuf17, spc17_phy_pc_w[8:1]};
       if (spc17_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 17, linebuf17);
          linebuf17 = "";
       end
    end else begin
       hitMadPrint17 = 0;
    end
  end
end


string linebuf18 = "";
logic hitMadPrint18 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc18_inst_done && ((spc18_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint18 = 1;
       linebuf18 = {linebuf18, spc18_phy_pc_w[8:1]};
       if (spc18_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 18, linebuf18);
          linebuf18 = "";
       end
    end else begin
       hitMadPrint18 = 0;
    end
  end
end


string linebuf19 = "";
logic hitMadPrint19 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc19_inst_done && ((spc19_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint19 = 1;
       linebuf19 = {linebuf19, spc19_phy_pc_w[8:1]};
       if (spc19_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 19, linebuf19);
          linebuf19 = "";
       end
    end else begin
       hitMadPrint19 = 0;
    end
  end
end


string linebuf20 = "";
logic hitMadPrint20 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc20_inst_done && ((spc20_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint20 = 1;
       linebuf20 = {linebuf20, spc20_phy_pc_w[8:1]};
       if (spc20_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 20, linebuf20);
          linebuf20 = "";
       end
    end else begin
       hitMadPrint20 = 0;
    end
  end
end


string linebuf21 = "";
logic hitMadPrint21 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc21_inst_done && ((spc21_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint21 = 1;
       linebuf21 = {linebuf21, spc21_phy_pc_w[8:1]};
       if (spc21_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 21, linebuf21);
          linebuf21 = "";
       end
    end else begin
       hitMadPrint21 = 0;
    end
  end
end


string linebuf22 = "";
logic hitMadPrint22 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc22_inst_done && ((spc22_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint22 = 1;
       linebuf22 = {linebuf22, spc22_phy_pc_w[8:1]};
       if (spc22_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 22, linebuf22);
          linebuf22 = "";
       end
    end else begin
       hitMadPrint22 = 0;
    end
  end
end


string linebuf23 = "";
logic hitMadPrint23 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc23_inst_done && ((spc23_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint23 = 1;
       linebuf23 = {linebuf23, spc23_phy_pc_w[8:1]};
       if (spc23_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 23, linebuf23);
          linebuf23 = "";
       end
    end else begin
       hitMadPrint23 = 0;
    end
  end
end


string linebuf24 = "";
logic hitMadPrint24 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc24_inst_done && ((spc24_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint24 = 1;
       linebuf24 = {linebuf24, spc24_phy_pc_w[8:1]};
       if (spc24_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 24, linebuf24);
          linebuf24 = "";
       end
    end else begin
       hitMadPrint24 = 0;
    end
  end
end


string linebuf25 = "";
logic hitMadPrint25 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc25_inst_done && ((spc25_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint25 = 1;
       linebuf25 = {linebuf25, spc25_phy_pc_w[8:1]};
       if (spc25_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 25, linebuf25);
          linebuf25 = "";
       end
    end else begin
       hitMadPrint25 = 0;
    end
  end
end


string linebuf26 = "";
logic hitMadPrint26 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc26_inst_done && ((spc26_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint26 = 1;
       linebuf26 = {linebuf26, spc26_phy_pc_w[8:1]};
       if (spc26_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 26, linebuf26);
          linebuf26 = "";
       end
    end else begin
       hitMadPrint26 = 0;
    end
  end
end


string linebuf27 = "";
logic hitMadPrint27 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc27_inst_done && ((spc27_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint27 = 1;
       linebuf27 = {linebuf27, spc27_phy_pc_w[8:1]};
       if (spc27_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 27, linebuf27);
          linebuf27 = "";
       end
    end else begin
       hitMadPrint27 = 0;
    end
  end
end


string linebuf28 = "";
logic hitMadPrint28 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc28_inst_done && ((spc28_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint28 = 1;
       linebuf28 = {linebuf28, spc28_phy_pc_w[8:1]};
       if (spc28_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 28, linebuf28);
          linebuf28 = "";
       end
    end else begin
       hitMadPrint28 = 0;
    end
  end
end


string linebuf29 = "";
logic hitMadPrint29 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc29_inst_done && ((spc29_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint29 = 1;
       linebuf29 = {linebuf29, spc29_phy_pc_w[8:1]};
       if (spc29_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 29, linebuf29);
          linebuf29 = "";
       end
    end else begin
       hitMadPrint29 = 0;
    end
  end
end


string linebuf30 = "";
logic hitMadPrint30 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc30_inst_done && ((spc30_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint30 = 1;
       linebuf30 = {linebuf30, spc30_phy_pc_w[8:1]};
       if (spc30_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 30, linebuf30);
          linebuf30 = "";
       end
    end else begin
       hitMadPrint30 = 0;
    end
  end
end


string linebuf31 = "";
logic hitMadPrint31 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc31_inst_done && ((spc31_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint31 = 1;
       linebuf31 = {linebuf31, spc31_phy_pc_w[8:1]};
       if (spc31_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 31, linebuf31);
          linebuf31 = "";
       end
    end else begin
       hitMadPrint31 = 0;
    end
  end
end


string linebuf32 = "";
logic hitMadPrint32 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc32_inst_done && ((spc32_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint32 = 1;
       linebuf32 = {linebuf32, spc32_phy_pc_w[8:1]};
       if (spc32_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 32, linebuf32);
          linebuf32 = "";
       end
    end else begin
       hitMadPrint32 = 0;
    end
  end
end


string linebuf33 = "";
logic hitMadPrint33 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc33_inst_done && ((spc33_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint33 = 1;
       linebuf33 = {linebuf33, spc33_phy_pc_w[8:1]};
       if (spc33_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 33, linebuf33);
          linebuf33 = "";
       end
    end else begin
       hitMadPrint33 = 0;
    end
  end
end


string linebuf34 = "";
logic hitMadPrint34 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc34_inst_done && ((spc34_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint34 = 1;
       linebuf34 = {linebuf34, spc34_phy_pc_w[8:1]};
       if (spc34_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 34, linebuf34);
          linebuf34 = "";
       end
    end else begin
       hitMadPrint34 = 0;
    end
  end
end


string linebuf35 = "";
logic hitMadPrint35 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc35_inst_done && ((spc35_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint35 = 1;
       linebuf35 = {linebuf35, spc35_phy_pc_w[8:1]};
       if (spc35_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 35, linebuf35);
          linebuf35 = "";
       end
    end else begin
       hitMadPrint35 = 0;
    end
  end
end


string linebuf36 = "";
logic hitMadPrint36 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc36_inst_done && ((spc36_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint36 = 1;
       linebuf36 = {linebuf36, spc36_phy_pc_w[8:1]};
       if (spc36_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 36, linebuf36);
          linebuf36 = "";
       end
    end else begin
       hitMadPrint36 = 0;
    end
  end
end


string linebuf37 = "";
logic hitMadPrint37 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc37_inst_done && ((spc37_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint37 = 1;
       linebuf37 = {linebuf37, spc37_phy_pc_w[8:1]};
       if (spc37_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 37, linebuf37);
          linebuf37 = "";
       end
    end else begin
       hitMadPrint37 = 0;
    end
  end
end


string linebuf38 = "";
logic hitMadPrint38 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc38_inst_done && ((spc38_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint38 = 1;
       linebuf38 = {linebuf38, spc38_phy_pc_w[8:1]};
       if (spc38_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 38, linebuf38);
          linebuf38 = "";
       end
    end else begin
       hitMadPrint38 = 0;
    end
  end
end


string linebuf39 = "";
logic hitMadPrint39 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc39_inst_done && ((spc39_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint39 = 1;
       linebuf39 = {linebuf39, spc39_phy_pc_w[8:1]};
       if (spc39_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 39, linebuf39);
          linebuf39 = "";
       end
    end else begin
       hitMadPrint39 = 0;
    end
  end
end


string linebuf40 = "";
logic hitMadPrint40 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc40_inst_done && ((spc40_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint40 = 1;
       linebuf40 = {linebuf40, spc40_phy_pc_w[8:1]};
       if (spc40_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 40, linebuf40);
          linebuf40 = "";
       end
    end else begin
       hitMadPrint40 = 0;
    end
  end
end


string linebuf41 = "";
logic hitMadPrint41 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc41_inst_done && ((spc41_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint41 = 1;
       linebuf41 = {linebuf41, spc41_phy_pc_w[8:1]};
       if (spc41_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 41, linebuf41);
          linebuf41 = "";
       end
    end else begin
       hitMadPrint41 = 0;
    end
  end
end


string linebuf42 = "";
logic hitMadPrint42 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc42_inst_done && ((spc42_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint42 = 1;
       linebuf42 = {linebuf42, spc42_phy_pc_w[8:1]};
       if (spc42_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 42, linebuf42);
          linebuf42 = "";
       end
    end else begin
       hitMadPrint42 = 0;
    end
  end
end


string linebuf43 = "";
logic hitMadPrint43 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc43_inst_done && ((spc43_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint43 = 1;
       linebuf43 = {linebuf43, spc43_phy_pc_w[8:1]};
       if (spc43_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 43, linebuf43);
          linebuf43 = "";
       end
    end else begin
       hitMadPrint43 = 0;
    end
  end
end


string linebuf44 = "";
logic hitMadPrint44 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc44_inst_done && ((spc44_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint44 = 1;
       linebuf44 = {linebuf44, spc44_phy_pc_w[8:1]};
       if (spc44_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 44, linebuf44);
          linebuf44 = "";
       end
    end else begin
       hitMadPrint44 = 0;
    end
  end
end


string linebuf45 = "";
logic hitMadPrint45 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc45_inst_done && ((spc45_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint45 = 1;
       linebuf45 = {linebuf45, spc45_phy_pc_w[8:1]};
       if (spc45_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 45, linebuf45);
          linebuf45 = "";
       end
    end else begin
       hitMadPrint45 = 0;
    end
  end
end


string linebuf46 = "";
logic hitMadPrint46 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc46_inst_done && ((spc46_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint46 = 1;
       linebuf46 = {linebuf46, spc46_phy_pc_w[8:1]};
       if (spc46_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 46, linebuf46);
          linebuf46 = "";
       end
    end else begin
       hitMadPrint46 = 0;
    end
  end
end


string linebuf47 = "";
logic hitMadPrint47 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc47_inst_done && ((spc47_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint47 = 1;
       linebuf47 = {linebuf47, spc47_phy_pc_w[8:1]};
       if (spc47_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 47, linebuf47);
          linebuf47 = "";
       end
    end else begin
       hitMadPrint47 = 0;
    end
  end
end


string linebuf48 = "";
logic hitMadPrint48 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc48_inst_done && ((spc48_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint48 = 1;
       linebuf48 = {linebuf48, spc48_phy_pc_w[8:1]};
       if (spc48_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 48, linebuf48);
          linebuf48 = "";
       end
    end else begin
       hitMadPrint48 = 0;
    end
  end
end


string linebuf49 = "";
logic hitMadPrint49 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc49_inst_done && ((spc49_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint49 = 1;
       linebuf49 = {linebuf49, spc49_phy_pc_w[8:1]};
       if (spc49_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 49, linebuf49);
          linebuf49 = "";
       end
    end else begin
       hitMadPrint49 = 0;
    end
  end
end


string linebuf50 = "";
logic hitMadPrint50 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc50_inst_done && ((spc50_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint50 = 1;
       linebuf50 = {linebuf50, spc50_phy_pc_w[8:1]};
       if (spc50_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 50, linebuf50);
          linebuf50 = "";
       end
    end else begin
       hitMadPrint50 = 0;
    end
  end
end


string linebuf51 = "";
logic hitMadPrint51 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc51_inst_done && ((spc51_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint51 = 1;
       linebuf51 = {linebuf51, spc51_phy_pc_w[8:1]};
       if (spc51_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 51, linebuf51);
          linebuf51 = "";
       end
    end else begin
       hitMadPrint51 = 0;
    end
  end
end


string linebuf52 = "";
logic hitMadPrint52 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc52_inst_done && ((spc52_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint52 = 1;
       linebuf52 = {linebuf52, spc52_phy_pc_w[8:1]};
       if (spc52_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 52, linebuf52);
          linebuf52 = "";
       end
    end else begin
       hitMadPrint52 = 0;
    end
  end
end


string linebuf53 = "";
logic hitMadPrint53 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc53_inst_done && ((spc53_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint53 = 1;
       linebuf53 = {linebuf53, spc53_phy_pc_w[8:1]};
       if (spc53_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 53, linebuf53);
          linebuf53 = "";
       end
    end else begin
       hitMadPrint53 = 0;
    end
  end
end


string linebuf54 = "";
logic hitMadPrint54 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc54_inst_done && ((spc54_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint54 = 1;
       linebuf54 = {linebuf54, spc54_phy_pc_w[8:1]};
       if (spc54_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 54, linebuf54);
          linebuf54 = "";
       end
    end else begin
       hitMadPrint54 = 0;
    end
  end
end


string linebuf55 = "";
logic hitMadPrint55 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc55_inst_done && ((spc55_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint55 = 1;
       linebuf55 = {linebuf55, spc55_phy_pc_w[8:1]};
       if (spc55_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 55, linebuf55);
          linebuf55 = "";
       end
    end else begin
       hitMadPrint55 = 0;
    end
  end
end


string linebuf56 = "";
logic hitMadPrint56 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc56_inst_done && ((spc56_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint56 = 1;
       linebuf56 = {linebuf56, spc56_phy_pc_w[8:1]};
       if (spc56_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 56, linebuf56);
          linebuf56 = "";
       end
    end else begin
       hitMadPrint56 = 0;
    end
  end
end


string linebuf57 = "";
logic hitMadPrint57 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc57_inst_done && ((spc57_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint57 = 1;
       linebuf57 = {linebuf57, spc57_phy_pc_w[8:1]};
       if (spc57_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 57, linebuf57);
          linebuf57 = "";
       end
    end else begin
       hitMadPrint57 = 0;
    end
  end
end


string linebuf58 = "";
logic hitMadPrint58 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc58_inst_done && ((spc58_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint58 = 1;
       linebuf58 = {linebuf58, spc58_phy_pc_w[8:1]};
       if (spc58_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 58, linebuf58);
          linebuf58 = "";
       end
    end else begin
       hitMadPrint58 = 0;
    end
  end
end


string linebuf59 = "";
logic hitMadPrint59 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc59_inst_done && ((spc59_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint59 = 1;
       linebuf59 = {linebuf59, spc59_phy_pc_w[8:1]};
       if (spc59_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 59, linebuf59);
          linebuf59 = "";
       end
    end else begin
       hitMadPrint59 = 0;
    end
  end
end


string linebuf60 = "";
logic hitMadPrint60 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc60_inst_done && ((spc60_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint60 = 1;
       linebuf60 = {linebuf60, spc60_phy_pc_w[8:1]};
       if (spc60_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 60, linebuf60);
          linebuf60 = "";
       end
    end else begin
       hitMadPrint60 = 0;
    end
  end
end


string linebuf61 = "";
logic hitMadPrint61 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc61_inst_done && ((spc61_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint61 = 1;
       linebuf61 = {linebuf61, spc61_phy_pc_w[8:1]};
       if (spc61_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 61, linebuf61);
          linebuf61 = "";
       end
    end else begin
       hitMadPrint61 = 0;
    end
  end
end


string linebuf62 = "";
logic hitMadPrint62 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc62_inst_done && ((spc62_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint62 = 1;
       linebuf62 = {linebuf62, spc62_phy_pc_w[8:1]};
       if (spc62_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 62, linebuf62);
          linebuf62 = "";
       end
    end else begin
       hitMadPrint62 = 0;
    end
  end
end


string linebuf63 = "";
logic hitMadPrint63 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc63_inst_done && ((spc63_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint63 = 1;
       linebuf63 = {linebuf63, spc63_phy_pc_w[8:1]};
       if (spc63_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 63, linebuf63);
          linebuf63 = "";
       end
    end else begin
       hitMadPrint63 = 0;
    end
  end
end


string linebuf64 = "";
logic hitMadPrint64 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc64_inst_done && ((spc64_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint64 = 1;
       linebuf64 = {linebuf64, spc64_phy_pc_w[8:1]};
       if (spc64_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 64, linebuf64);
          linebuf64 = "";
       end
    end else begin
       hitMadPrint64 = 0;
    end
  end
end


string linebuf65 = "";
logic hitMadPrint65 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc65_inst_done && ((spc65_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint65 = 1;
       linebuf65 = {linebuf65, spc65_phy_pc_w[8:1]};
       if (spc65_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 65, linebuf65);
          linebuf65 = "";
       end
    end else begin
       hitMadPrint65 = 0;
    end
  end
end


string linebuf66 = "";
logic hitMadPrint66 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc66_inst_done && ((spc66_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint66 = 1;
       linebuf66 = {linebuf66, spc66_phy_pc_w[8:1]};
       if (spc66_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 66, linebuf66);
          linebuf66 = "";
       end
    end else begin
       hitMadPrint66 = 0;
    end
  end
end


string linebuf67 = "";
logic hitMadPrint67 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc67_inst_done && ((spc67_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint67 = 1;
       linebuf67 = {linebuf67, spc67_phy_pc_w[8:1]};
       if (spc67_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 67, linebuf67);
          linebuf67 = "";
       end
    end else begin
       hitMadPrint67 = 0;
    end
  end
end


string linebuf68 = "";
logic hitMadPrint68 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc68_inst_done && ((spc68_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint68 = 1;
       linebuf68 = {linebuf68, spc68_phy_pc_w[8:1]};
       if (spc68_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 68, linebuf68);
          linebuf68 = "";
       end
    end else begin
       hitMadPrint68 = 0;
    end
  end
end


string linebuf69 = "";
logic hitMadPrint69 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc69_inst_done && ((spc69_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint69 = 1;
       linebuf69 = {linebuf69, spc69_phy_pc_w[8:1]};
       if (spc69_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 69, linebuf69);
          linebuf69 = "";
       end
    end else begin
       hitMadPrint69 = 0;
    end
  end
end


string linebuf70 = "";
logic hitMadPrint70 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc70_inst_done && ((spc70_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint70 = 1;
       linebuf70 = {linebuf70, spc70_phy_pc_w[8:1]};
       if (spc70_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 70, linebuf70);
          linebuf70 = "";
       end
    end else begin
       hitMadPrint70 = 0;
    end
  end
end


string linebuf71 = "";
logic hitMadPrint71 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc71_inst_done && ((spc71_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint71 = 1;
       linebuf71 = {linebuf71, spc71_phy_pc_w[8:1]};
       if (spc71_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 71, linebuf71);
          linebuf71 = "";
       end
    end else begin
       hitMadPrint71 = 0;
    end
  end
end


string linebuf72 = "";
logic hitMadPrint72 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc72_inst_done && ((spc72_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint72 = 1;
       linebuf72 = {linebuf72, spc72_phy_pc_w[8:1]};
       if (spc72_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 72, linebuf72);
          linebuf72 = "";
       end
    end else begin
       hitMadPrint72 = 0;
    end
  end
end


string linebuf73 = "";
logic hitMadPrint73 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc73_inst_done && ((spc73_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint73 = 1;
       linebuf73 = {linebuf73, spc73_phy_pc_w[8:1]};
       if (spc73_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 73, linebuf73);
          linebuf73 = "";
       end
    end else begin
       hitMadPrint73 = 0;
    end
  end
end


string linebuf74 = "";
logic hitMadPrint74 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc74_inst_done && ((spc74_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint74 = 1;
       linebuf74 = {linebuf74, spc74_phy_pc_w[8:1]};
       if (spc74_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 74, linebuf74);
          linebuf74 = "";
       end
    end else begin
       hitMadPrint74 = 0;
    end
  end
end


string linebuf75 = "";
logic hitMadPrint75 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc75_inst_done && ((spc75_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint75 = 1;
       linebuf75 = {linebuf75, spc75_phy_pc_w[8:1]};
       if (spc75_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 75, linebuf75);
          linebuf75 = "";
       end
    end else begin
       hitMadPrint75 = 0;
    end
  end
end


string linebuf76 = "";
logic hitMadPrint76 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc76_inst_done && ((spc76_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint76 = 1;
       linebuf76 = {linebuf76, spc76_phy_pc_w[8:1]};
       if (spc76_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 76, linebuf76);
          linebuf76 = "";
       end
    end else begin
       hitMadPrint76 = 0;
    end
  end
end


string linebuf77 = "";
logic hitMadPrint77 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc77_inst_done && ((spc77_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint77 = 1;
       linebuf77 = {linebuf77, spc77_phy_pc_w[8:1]};
       if (spc77_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 77, linebuf77);
          linebuf77 = "";
       end
    end else begin
       hitMadPrint77 = 0;
    end
  end
end


string linebuf78 = "";
logic hitMadPrint78 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc78_inst_done && ((spc78_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint78 = 1;
       linebuf78 = {linebuf78, spc78_phy_pc_w[8:1]};
       if (spc78_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 78, linebuf78);
          linebuf78 = "";
       end
    end else begin
       hitMadPrint78 = 0;
    end
  end
end


string linebuf79 = "";
logic hitMadPrint79 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc79_inst_done && ((spc79_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint79 = 1;
       linebuf79 = {linebuf79, spc79_phy_pc_w[8:1]};
       if (spc79_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 79, linebuf79);
          linebuf79 = "";
       end
    end else begin
       hitMadPrint79 = 0;
    end
  end
end


string linebuf80 = "";
logic hitMadPrint80 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc80_inst_done && ((spc80_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint80 = 1;
       linebuf80 = {linebuf80, spc80_phy_pc_w[8:1]};
       if (spc80_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 80, linebuf80);
          linebuf80 = "";
       end
    end else begin
       hitMadPrint80 = 0;
    end
  end
end


string linebuf81 = "";
logic hitMadPrint81 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc81_inst_done && ((spc81_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint81 = 1;
       linebuf81 = {linebuf81, spc81_phy_pc_w[8:1]};
       if (spc81_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 81, linebuf81);
          linebuf81 = "";
       end
    end else begin
       hitMadPrint81 = 0;
    end
  end
end


string linebuf82 = "";
logic hitMadPrint82 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc82_inst_done && ((spc82_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint82 = 1;
       linebuf82 = {linebuf82, spc82_phy_pc_w[8:1]};
       if (spc82_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 82, linebuf82);
          linebuf82 = "";
       end
    end else begin
       hitMadPrint82 = 0;
    end
  end
end


string linebuf83 = "";
logic hitMadPrint83 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc83_inst_done && ((spc83_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint83 = 1;
       linebuf83 = {linebuf83, spc83_phy_pc_w[8:1]};
       if (spc83_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 83, linebuf83);
          linebuf83 = "";
       end
    end else begin
       hitMadPrint83 = 0;
    end
  end
end


string linebuf84 = "";
logic hitMadPrint84 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc84_inst_done && ((spc84_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint84 = 1;
       linebuf84 = {linebuf84, spc84_phy_pc_w[8:1]};
       if (spc84_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 84, linebuf84);
          linebuf84 = "";
       end
    end else begin
       hitMadPrint84 = 0;
    end
  end
end


string linebuf85 = "";
logic hitMadPrint85 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc85_inst_done && ((spc85_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint85 = 1;
       linebuf85 = {linebuf85, spc85_phy_pc_w[8:1]};
       if (spc85_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 85, linebuf85);
          linebuf85 = "";
       end
    end else begin
       hitMadPrint85 = 0;
    end
  end
end


string linebuf86 = "";
logic hitMadPrint86 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc86_inst_done && ((spc86_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint86 = 1;
       linebuf86 = {linebuf86, spc86_phy_pc_w[8:1]};
       if (spc86_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 86, linebuf86);
          linebuf86 = "";
       end
    end else begin
       hitMadPrint86 = 0;
    end
  end
end


string linebuf87 = "";
logic hitMadPrint87 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc87_inst_done && ((spc87_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint87 = 1;
       linebuf87 = {linebuf87, spc87_phy_pc_w[8:1]};
       if (spc87_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 87, linebuf87);
          linebuf87 = "";
       end
    end else begin
       hitMadPrint87 = 0;
    end
  end
end


string linebuf88 = "";
logic hitMadPrint88 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc88_inst_done && ((spc88_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint88 = 1;
       linebuf88 = {linebuf88, spc88_phy_pc_w[8:1]};
       if (spc88_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 88, linebuf88);
          linebuf88 = "";
       end
    end else begin
       hitMadPrint88 = 0;
    end
  end
end


string linebuf89 = "";
logic hitMadPrint89 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc89_inst_done && ((spc89_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint89 = 1;
       linebuf89 = {linebuf89, spc89_phy_pc_w[8:1]};
       if (spc89_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 89, linebuf89);
          linebuf89 = "";
       end
    end else begin
       hitMadPrint89 = 0;
    end
  end
end


string linebuf90 = "";
logic hitMadPrint90 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc90_inst_done && ((spc90_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint90 = 1;
       linebuf90 = {linebuf90, spc90_phy_pc_w[8:1]};
       if (spc90_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 90, linebuf90);
          linebuf90 = "";
       end
    end else begin
       hitMadPrint90 = 0;
    end
  end
end


string linebuf91 = "";
logic hitMadPrint91 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc91_inst_done && ((spc91_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint91 = 1;
       linebuf91 = {linebuf91, spc91_phy_pc_w[8:1]};
       if (spc91_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 91, linebuf91);
          linebuf91 = "";
       end
    end else begin
       hitMadPrint91 = 0;
    end
  end
end


string linebuf92 = "";
logic hitMadPrint92 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc92_inst_done && ((spc92_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint92 = 1;
       linebuf92 = {linebuf92, spc92_phy_pc_w[8:1]};
       if (spc92_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 92, linebuf92);
          linebuf92 = "";
       end
    end else begin
       hitMadPrint92 = 0;
    end
  end
end


string linebuf93 = "";
logic hitMadPrint93 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc93_inst_done && ((spc93_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint93 = 1;
       linebuf93 = {linebuf93, spc93_phy_pc_w[8:1]};
       if (spc93_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 93, linebuf93);
          linebuf93 = "";
       end
    end else begin
       hitMadPrint93 = 0;
    end
  end
end


string linebuf94 = "";
logic hitMadPrint94 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc94_inst_done && ((spc94_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint94 = 1;
       linebuf94 = {linebuf94, spc94_phy_pc_w[8:1]};
       if (spc94_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 94, linebuf94);
          linebuf94 = "";
       end
    end else begin
       hitMadPrint94 = 0;
    end
  end
end


string linebuf95 = "";
logic hitMadPrint95 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc95_inst_done && ((spc95_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint95 = 1;
       linebuf95 = {linebuf95, spc95_phy_pc_w[8:1]};
       if (spc95_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 95, linebuf95);
          linebuf95 = "";
       end
    end else begin
       hitMadPrint95 = 0;
    end
  end
end


string linebuf96 = "";
logic hitMadPrint96 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc96_inst_done && ((spc96_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint96 = 1;
       linebuf96 = {linebuf96, spc96_phy_pc_w[8:1]};
       if (spc96_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 96, linebuf96);
          linebuf96 = "";
       end
    end else begin
       hitMadPrint96 = 0;
    end
  end
end


string linebuf97 = "";
logic hitMadPrint97 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc97_inst_done && ((spc97_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint97 = 1;
       linebuf97 = {linebuf97, spc97_phy_pc_w[8:1]};
       if (spc97_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 97, linebuf97);
          linebuf97 = "";
       end
    end else begin
       hitMadPrint97 = 0;
    end
  end
end


string linebuf98 = "";
logic hitMadPrint98 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc98_inst_done && ((spc98_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint98 = 1;
       linebuf98 = {linebuf98, spc98_phy_pc_w[8:1]};
       if (spc98_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 98, linebuf98);
          linebuf98 = "";
       end
    end else begin
       hitMadPrint98 = 0;
    end
  end
end


string linebuf99 = "";
logic hitMadPrint99 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc99_inst_done && ((spc99_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint99 = 1;
       linebuf99 = {linebuf99, spc99_phy_pc_w[8:1]};
       if (spc99_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 99, linebuf99);
          linebuf99 = "";
       end
    end else begin
       hitMadPrint99 = 0;
    end
  end
end


string linebuf100 = "";
logic hitMadPrint100 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc100_inst_done && ((spc100_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint100 = 1;
       linebuf100 = {linebuf100, spc100_phy_pc_w[8:1]};
       if (spc100_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 100, linebuf100);
          linebuf100 = "";
       end
    end else begin
       hitMadPrint100 = 0;
    end
  end
end


string linebuf101 = "";
logic hitMadPrint101 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc101_inst_done && ((spc101_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint101 = 1;
       linebuf101 = {linebuf101, spc101_phy_pc_w[8:1]};
       if (spc101_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 101, linebuf101);
          linebuf101 = "";
       end
    end else begin
       hitMadPrint101 = 0;
    end
  end
end


string linebuf102 = "";
logic hitMadPrint102 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc102_inst_done && ((spc102_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint102 = 1;
       linebuf102 = {linebuf102, spc102_phy_pc_w[8:1]};
       if (spc102_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 102, linebuf102);
          linebuf102 = "";
       end
    end else begin
       hitMadPrint102 = 0;
    end
  end
end


string linebuf103 = "";
logic hitMadPrint103 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc103_inst_done && ((spc103_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint103 = 1;
       linebuf103 = {linebuf103, spc103_phy_pc_w[8:1]};
       if (spc103_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 103, linebuf103);
          linebuf103 = "";
       end
    end else begin
       hitMadPrint103 = 0;
    end
  end
end


string linebuf104 = "";
logic hitMadPrint104 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc104_inst_done && ((spc104_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint104 = 1;
       linebuf104 = {linebuf104, spc104_phy_pc_w[8:1]};
       if (spc104_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 104, linebuf104);
          linebuf104 = "";
       end
    end else begin
       hitMadPrint104 = 0;
    end
  end
end


string linebuf105 = "";
logic hitMadPrint105 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc105_inst_done && ((spc105_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint105 = 1;
       linebuf105 = {linebuf105, spc105_phy_pc_w[8:1]};
       if (spc105_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 105, linebuf105);
          linebuf105 = "";
       end
    end else begin
       hitMadPrint105 = 0;
    end
  end
end


string linebuf106 = "";
logic hitMadPrint106 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc106_inst_done && ((spc106_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint106 = 1;
       linebuf106 = {linebuf106, spc106_phy_pc_w[8:1]};
       if (spc106_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 106, linebuf106);
          linebuf106 = "";
       end
    end else begin
       hitMadPrint106 = 0;
    end
  end
end


string linebuf107 = "";
logic hitMadPrint107 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc107_inst_done && ((spc107_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint107 = 1;
       linebuf107 = {linebuf107, spc107_phy_pc_w[8:1]};
       if (spc107_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 107, linebuf107);
          linebuf107 = "";
       end
    end else begin
       hitMadPrint107 = 0;
    end
  end
end


string linebuf108 = "";
logic hitMadPrint108 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc108_inst_done && ((spc108_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint108 = 1;
       linebuf108 = {linebuf108, spc108_phy_pc_w[8:1]};
       if (spc108_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 108, linebuf108);
          linebuf108 = "";
       end
    end else begin
       hitMadPrint108 = 0;
    end
  end
end


string linebuf109 = "";
logic hitMadPrint109 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc109_inst_done && ((spc109_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint109 = 1;
       linebuf109 = {linebuf109, spc109_phy_pc_w[8:1]};
       if (spc109_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 109, linebuf109);
          linebuf109 = "";
       end
    end else begin
       hitMadPrint109 = 0;
    end
  end
end


string linebuf110 = "";
logic hitMadPrint110 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc110_inst_done && ((spc110_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint110 = 1;
       linebuf110 = {linebuf110, spc110_phy_pc_w[8:1]};
       if (spc110_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 110, linebuf110);
          linebuf110 = "";
       end
    end else begin
       hitMadPrint110 = 0;
    end
  end
end


string linebuf111 = "";
logic hitMadPrint111 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc111_inst_done && ((spc111_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint111 = 1;
       linebuf111 = {linebuf111, spc111_phy_pc_w[8:1]};
       if (spc111_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 111, linebuf111);
          linebuf111 = "";
       end
    end else begin
       hitMadPrint111 = 0;
    end
  end
end


string linebuf112 = "";
logic hitMadPrint112 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc112_inst_done && ((spc112_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint112 = 1;
       linebuf112 = {linebuf112, spc112_phy_pc_w[8:1]};
       if (spc112_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 112, linebuf112);
          linebuf112 = "";
       end
    end else begin
       hitMadPrint112 = 0;
    end
  end
end


string linebuf113 = "";
logic hitMadPrint113 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc113_inst_done && ((spc113_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint113 = 1;
       linebuf113 = {linebuf113, spc113_phy_pc_w[8:1]};
       if (spc113_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 113, linebuf113);
          linebuf113 = "";
       end
    end else begin
       hitMadPrint113 = 0;
    end
  end
end


string linebuf114 = "";
logic hitMadPrint114 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc114_inst_done && ((spc114_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint114 = 1;
       linebuf114 = {linebuf114, spc114_phy_pc_w[8:1]};
       if (spc114_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 114, linebuf114);
          linebuf114 = "";
       end
    end else begin
       hitMadPrint114 = 0;
    end
  end
end


string linebuf115 = "";
logic hitMadPrint115 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc115_inst_done && ((spc115_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint115 = 1;
       linebuf115 = {linebuf115, spc115_phy_pc_w[8:1]};
       if (spc115_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 115, linebuf115);
          linebuf115 = "";
       end
    end else begin
       hitMadPrint115 = 0;
    end
  end
end


string linebuf116 = "";
logic hitMadPrint116 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc116_inst_done && ((spc116_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint116 = 1;
       linebuf116 = {linebuf116, spc116_phy_pc_w[8:1]};
       if (spc116_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 116, linebuf116);
          linebuf116 = "";
       end
    end else begin
       hitMadPrint116 = 0;
    end
  end
end


string linebuf117 = "";
logic hitMadPrint117 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc117_inst_done && ((spc117_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint117 = 1;
       linebuf117 = {linebuf117, spc117_phy_pc_w[8:1]};
       if (spc117_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 117, linebuf117);
          linebuf117 = "";
       end
    end else begin
       hitMadPrint117 = 0;
    end
  end
end


string linebuf118 = "";
logic hitMadPrint118 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc118_inst_done && ((spc118_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint118 = 1;
       linebuf118 = {linebuf118, spc118_phy_pc_w[8:1]};
       if (spc118_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 118, linebuf118);
          linebuf118 = "";
       end
    end else begin
       hitMadPrint118 = 0;
    end
  end
end


string linebuf119 = "";
logic hitMadPrint119 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc119_inst_done && ((spc119_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint119 = 1;
       linebuf119 = {linebuf119, spc119_phy_pc_w[8:1]};
       if (spc119_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 119, linebuf119);
          linebuf119 = "";
       end
    end else begin
       hitMadPrint119 = 0;
    end
  end
end


string linebuf120 = "";
logic hitMadPrint120 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc120_inst_done && ((spc120_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint120 = 1;
       linebuf120 = {linebuf120, spc120_phy_pc_w[8:1]};
       if (spc120_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 120, linebuf120);
          linebuf120 = "";
       end
    end else begin
       hitMadPrint120 = 0;
    end
  end
end


string linebuf121 = "";
logic hitMadPrint121 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc121_inst_done && ((spc121_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint121 = 1;
       linebuf121 = {linebuf121, spc121_phy_pc_w[8:1]};
       if (spc121_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 121, linebuf121);
          linebuf121 = "";
       end
    end else begin
       hitMadPrint121 = 0;
    end
  end
end


string linebuf122 = "";
logic hitMadPrint122 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc122_inst_done && ((spc122_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint122 = 1;
       linebuf122 = {linebuf122, spc122_phy_pc_w[8:1]};
       if (spc122_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 122, linebuf122);
          linebuf122 = "";
       end
    end else begin
       hitMadPrint122 = 0;
    end
  end
end


string linebuf123 = "";
logic hitMadPrint123 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc123_inst_done && ((spc123_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint123 = 1;
       linebuf123 = {linebuf123, spc123_phy_pc_w[8:1]};
       if (spc123_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 123, linebuf123);
          linebuf123 = "";
       end
    end else begin
       hitMadPrint123 = 0;
    end
  end
end


string linebuf124 = "";
logic hitMadPrint124 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc124_inst_done && ((spc124_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint124 = 1;
       linebuf124 = {linebuf124, spc124_phy_pc_w[8:1]};
       if (spc124_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 124, linebuf124);
          linebuf124 = "";
       end
    end else begin
       hitMadPrint124 = 0;
    end
  end
end


string linebuf125 = "";
logic hitMadPrint125 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc125_inst_done && ((spc125_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint125 = 1;
       linebuf125 = {linebuf125, spc125_phy_pc_w[8:1]};
       if (spc125_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 125, linebuf125);
          linebuf125 = "";
       end
    end else begin
       hitMadPrint125 = 0;
    end
  end
end


string linebuf126 = "";
logic hitMadPrint126 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc126_inst_done && ((spc126_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint126 = 1;
       linebuf126 = {linebuf126, spc126_phy_pc_w[8:1]};
       if (spc126_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 126, linebuf126);
          linebuf126 = "";
       end
    end else begin
       hitMadPrint126 = 0;
    end
  end
end


string linebuf127 = "";
logic hitMadPrint127 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc127_inst_done && ((spc127_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint127 = 1;
       linebuf127 = {linebuf127, spc127_phy_pc_w[8:1]};
       if (spc127_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 127, linebuf127);
          linebuf127 = "";
       end
    end else begin
       hitMadPrint127 = 0;
    end
  end
end


string linebuf128 = "";
logic hitMadPrint128 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc128_inst_done && ((spc128_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint128 = 1;
       linebuf128 = {linebuf128, spc128_phy_pc_w[8:1]};
       if (spc128_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 128, linebuf128);
          linebuf128 = "";
       end
    end else begin
       hitMadPrint128 = 0;
    end
  end
end


string linebuf129 = "";
logic hitMadPrint129 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc129_inst_done && ((spc129_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint129 = 1;
       linebuf129 = {linebuf129, spc129_phy_pc_w[8:1]};
       if (spc129_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 129, linebuf129);
          linebuf129 = "";
       end
    end else begin
       hitMadPrint129 = 0;
    end
  end
end


string linebuf130 = "";
logic hitMadPrint130 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc130_inst_done && ((spc130_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint130 = 1;
       linebuf130 = {linebuf130, spc130_phy_pc_w[8:1]};
       if (spc130_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 130, linebuf130);
          linebuf130 = "";
       end
    end else begin
       hitMadPrint130 = 0;
    end
  end
end


string linebuf131 = "";
logic hitMadPrint131 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc131_inst_done && ((spc131_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint131 = 1;
       linebuf131 = {linebuf131, spc131_phy_pc_w[8:1]};
       if (spc131_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 131, linebuf131);
          linebuf131 = "";
       end
    end else begin
       hitMadPrint131 = 0;
    end
  end
end


string linebuf132 = "";
logic hitMadPrint132 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc132_inst_done && ((spc132_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint132 = 1;
       linebuf132 = {linebuf132, spc132_phy_pc_w[8:1]};
       if (spc132_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 132, linebuf132);
          linebuf132 = "";
       end
    end else begin
       hitMadPrint132 = 0;
    end
  end
end


string linebuf133 = "";
logic hitMadPrint133 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc133_inst_done && ((spc133_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint133 = 1;
       linebuf133 = {linebuf133, spc133_phy_pc_w[8:1]};
       if (spc133_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 133, linebuf133);
          linebuf133 = "";
       end
    end else begin
       hitMadPrint133 = 0;
    end
  end
end


string linebuf134 = "";
logic hitMadPrint134 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc134_inst_done && ((spc134_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint134 = 1;
       linebuf134 = {linebuf134, spc134_phy_pc_w[8:1]};
       if (spc134_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 134, linebuf134);
          linebuf134 = "";
       end
    end else begin
       hitMadPrint134 = 0;
    end
  end
end


string linebuf135 = "";
logic hitMadPrint135 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc135_inst_done && ((spc135_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint135 = 1;
       linebuf135 = {linebuf135, spc135_phy_pc_w[8:1]};
       if (spc135_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 135, linebuf135);
          linebuf135 = "";
       end
    end else begin
       hitMadPrint135 = 0;
    end
  end
end


string linebuf136 = "";
logic hitMadPrint136 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc136_inst_done && ((spc136_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint136 = 1;
       linebuf136 = {linebuf136, spc136_phy_pc_w[8:1]};
       if (spc136_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 136, linebuf136);
          linebuf136 = "";
       end
    end else begin
       hitMadPrint136 = 0;
    end
  end
end


string linebuf137 = "";
logic hitMadPrint137 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc137_inst_done && ((spc137_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint137 = 1;
       linebuf137 = {linebuf137, spc137_phy_pc_w[8:1]};
       if (spc137_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 137, linebuf137);
          linebuf137 = "";
       end
    end else begin
       hitMadPrint137 = 0;
    end
  end
end


string linebuf138 = "";
logic hitMadPrint138 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc138_inst_done && ((spc138_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint138 = 1;
       linebuf138 = {linebuf138, spc138_phy_pc_w[8:1]};
       if (spc138_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 138, linebuf138);
          linebuf138 = "";
       end
    end else begin
       hitMadPrint138 = 0;
    end
  end
end


string linebuf139 = "";
logic hitMadPrint139 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc139_inst_done && ((spc139_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint139 = 1;
       linebuf139 = {linebuf139, spc139_phy_pc_w[8:1]};
       if (spc139_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 139, linebuf139);
          linebuf139 = "";
       end
    end else begin
       hitMadPrint139 = 0;
    end
  end
end


string linebuf140 = "";
logic hitMadPrint140 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc140_inst_done && ((spc140_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint140 = 1;
       linebuf140 = {linebuf140, spc140_phy_pc_w[8:1]};
       if (spc140_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 140, linebuf140);
          linebuf140 = "";
       end
    end else begin
       hitMadPrint140 = 0;
    end
  end
end


string linebuf141 = "";
logic hitMadPrint141 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc141_inst_done && ((spc141_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint141 = 1;
       linebuf141 = {linebuf141, spc141_phy_pc_w[8:1]};
       if (spc141_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 141, linebuf141);
          linebuf141 = "";
       end
    end else begin
       hitMadPrint141 = 0;
    end
  end
end


string linebuf142 = "";
logic hitMadPrint142 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc142_inst_done && ((spc142_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint142 = 1;
       linebuf142 = {linebuf142, spc142_phy_pc_w[8:1]};
       if (spc142_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 142, linebuf142);
          linebuf142 = "";
       end
    end else begin
       hitMadPrint142 = 0;
    end
  end
end


string linebuf143 = "";
logic hitMadPrint143 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc143_inst_done && ((spc143_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint143 = 1;
       linebuf143 = {linebuf143, spc143_phy_pc_w[8:1]};
       if (spc143_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 143, linebuf143);
          linebuf143 = "";
       end
    end else begin
       hitMadPrint143 = 0;
    end
  end
end


string linebuf144 = "";
logic hitMadPrint144 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc144_inst_done && ((spc144_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint144 = 1;
       linebuf144 = {linebuf144, spc144_phy_pc_w[8:1]};
       if (spc144_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 144, linebuf144);
          linebuf144 = "";
       end
    end else begin
       hitMadPrint144 = 0;
    end
  end
end


string linebuf145 = "";
logic hitMadPrint145 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc145_inst_done && ((spc145_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint145 = 1;
       linebuf145 = {linebuf145, spc145_phy_pc_w[8:1]};
       if (spc145_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 145, linebuf145);
          linebuf145 = "";
       end
    end else begin
       hitMadPrint145 = 0;
    end
  end
end


string linebuf146 = "";
logic hitMadPrint146 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc146_inst_done && ((spc146_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint146 = 1;
       linebuf146 = {linebuf146, spc146_phy_pc_w[8:1]};
       if (spc146_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 146, linebuf146);
          linebuf146 = "";
       end
    end else begin
       hitMadPrint146 = 0;
    end
  end
end


string linebuf147 = "";
logic hitMadPrint147 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc147_inst_done && ((spc147_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint147 = 1;
       linebuf147 = {linebuf147, spc147_phy_pc_w[8:1]};
       if (spc147_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 147, linebuf147);
          linebuf147 = "";
       end
    end else begin
       hitMadPrint147 = 0;
    end
  end
end


string linebuf148 = "";
logic hitMadPrint148 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc148_inst_done && ((spc148_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint148 = 1;
       linebuf148 = {linebuf148, spc148_phy_pc_w[8:1]};
       if (spc148_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 148, linebuf148);
          linebuf148 = "";
       end
    end else begin
       hitMadPrint148 = 0;
    end
  end
end


string linebuf149 = "";
logic hitMadPrint149 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc149_inst_done && ((spc149_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint149 = 1;
       linebuf149 = {linebuf149, spc149_phy_pc_w[8:1]};
       if (spc149_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 149, linebuf149);
          linebuf149 = "";
       end
    end else begin
       hitMadPrint149 = 0;
    end
  end
end


string linebuf150 = "";
logic hitMadPrint150 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc150_inst_done && ((spc150_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint150 = 1;
       linebuf150 = {linebuf150, spc150_phy_pc_w[8:1]};
       if (spc150_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 150, linebuf150);
          linebuf150 = "";
       end
    end else begin
       hitMadPrint150 = 0;
    end
  end
end


string linebuf151 = "";
logic hitMadPrint151 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc151_inst_done && ((spc151_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint151 = 1;
       linebuf151 = {linebuf151, spc151_phy_pc_w[8:1]};
       if (spc151_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 151, linebuf151);
          linebuf151 = "";
       end
    end else begin
       hitMadPrint151 = 0;
    end
  end
end


string linebuf152 = "";
logic hitMadPrint152 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc152_inst_done && ((spc152_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint152 = 1;
       linebuf152 = {linebuf152, spc152_phy_pc_w[8:1]};
       if (spc152_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 152, linebuf152);
          linebuf152 = "";
       end
    end else begin
       hitMadPrint152 = 0;
    end
  end
end


string linebuf153 = "";
logic hitMadPrint153 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc153_inst_done && ((spc153_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint153 = 1;
       linebuf153 = {linebuf153, spc153_phy_pc_w[8:1]};
       if (spc153_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 153, linebuf153);
          linebuf153 = "";
       end
    end else begin
       hitMadPrint153 = 0;
    end
  end
end


string linebuf154 = "";
logic hitMadPrint154 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc154_inst_done && ((spc154_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint154 = 1;
       linebuf154 = {linebuf154, spc154_phy_pc_w[8:1]};
       if (spc154_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 154, linebuf154);
          linebuf154 = "";
       end
    end else begin
       hitMadPrint154 = 0;
    end
  end
end


string linebuf155 = "";
logic hitMadPrint155 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc155_inst_done && ((spc155_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint155 = 1;
       linebuf155 = {linebuf155, spc155_phy_pc_w[8:1]};
       if (spc155_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 155, linebuf155);
          linebuf155 = "";
       end
    end else begin
       hitMadPrint155 = 0;
    end
  end
end


string linebuf156 = "";
logic hitMadPrint156 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc156_inst_done && ((spc156_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint156 = 1;
       linebuf156 = {linebuf156, spc156_phy_pc_w[8:1]};
       if (spc156_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 156, linebuf156);
          linebuf156 = "";
       end
    end else begin
       hitMadPrint156 = 0;
    end
  end
end


string linebuf157 = "";
logic hitMadPrint157 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc157_inst_done && ((spc157_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint157 = 1;
       linebuf157 = {linebuf157, spc157_phy_pc_w[8:1]};
       if (spc157_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 157, linebuf157);
          linebuf157 = "";
       end
    end else begin
       hitMadPrint157 = 0;
    end
  end
end


string linebuf158 = "";
logic hitMadPrint158 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc158_inst_done && ((spc158_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint158 = 1;
       linebuf158 = {linebuf158, spc158_phy_pc_w[8:1]};
       if (spc158_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 158, linebuf158);
          linebuf158 = "";
       end
    end else begin
       hitMadPrint158 = 0;
    end
  end
end


string linebuf159 = "";
logic hitMadPrint159 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc159_inst_done && ((spc159_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint159 = 1;
       linebuf159 = {linebuf159, spc159_phy_pc_w[8:1]};
       if (spc159_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 159, linebuf159);
          linebuf159 = "";
       end
    end else begin
       hitMadPrint159 = 0;
    end
  end
end


string linebuf160 = "";
logic hitMadPrint160 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc160_inst_done && ((spc160_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint160 = 1;
       linebuf160 = {linebuf160, spc160_phy_pc_w[8:1]};
       if (spc160_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 160, linebuf160);
          linebuf160 = "";
       end
    end else begin
       hitMadPrint160 = 0;
    end
  end
end


string linebuf161 = "";
logic hitMadPrint161 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc161_inst_done && ((spc161_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint161 = 1;
       linebuf161 = {linebuf161, spc161_phy_pc_w[8:1]};
       if (spc161_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 161, linebuf161);
          linebuf161 = "";
       end
    end else begin
       hitMadPrint161 = 0;
    end
  end
end


string linebuf162 = "";
logic hitMadPrint162 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc162_inst_done && ((spc162_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint162 = 1;
       linebuf162 = {linebuf162, spc162_phy_pc_w[8:1]};
       if (spc162_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 162, linebuf162);
          linebuf162 = "";
       end
    end else begin
       hitMadPrint162 = 0;
    end
  end
end


string linebuf163 = "";
logic hitMadPrint163 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc163_inst_done && ((spc163_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint163 = 1;
       linebuf163 = {linebuf163, spc163_phy_pc_w[8:1]};
       if (spc163_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 163, linebuf163);
          linebuf163 = "";
       end
    end else begin
       hitMadPrint163 = 0;
    end
  end
end


string linebuf164 = "";
logic hitMadPrint164 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc164_inst_done && ((spc164_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint164 = 1;
       linebuf164 = {linebuf164, spc164_phy_pc_w[8:1]};
       if (spc164_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 164, linebuf164);
          linebuf164 = "";
       end
    end else begin
       hitMadPrint164 = 0;
    end
  end
end


string linebuf165 = "";
logic hitMadPrint165 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc165_inst_done && ((spc165_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint165 = 1;
       linebuf165 = {linebuf165, spc165_phy_pc_w[8:1]};
       if (spc165_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 165, linebuf165);
          linebuf165 = "";
       end
    end else begin
       hitMadPrint165 = 0;
    end
  end
end


string linebuf166 = "";
logic hitMadPrint166 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc166_inst_done && ((spc166_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint166 = 1;
       linebuf166 = {linebuf166, spc166_phy_pc_w[8:1]};
       if (spc166_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 166, linebuf166);
          linebuf166 = "";
       end
    end else begin
       hitMadPrint166 = 0;
    end
  end
end


string linebuf167 = "";
logic hitMadPrint167 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc167_inst_done && ((spc167_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint167 = 1;
       linebuf167 = {linebuf167, spc167_phy_pc_w[8:1]};
       if (spc167_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 167, linebuf167);
          linebuf167 = "";
       end
    end else begin
       hitMadPrint167 = 0;
    end
  end
end


string linebuf168 = "";
logic hitMadPrint168 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc168_inst_done && ((spc168_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint168 = 1;
       linebuf168 = {linebuf168, spc168_phy_pc_w[8:1]};
       if (spc168_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 168, linebuf168);
          linebuf168 = "";
       end
    end else begin
       hitMadPrint168 = 0;
    end
  end
end


string linebuf169 = "";
logic hitMadPrint169 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc169_inst_done && ((spc169_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint169 = 1;
       linebuf169 = {linebuf169, spc169_phy_pc_w[8:1]};
       if (spc169_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 169, linebuf169);
          linebuf169 = "";
       end
    end else begin
       hitMadPrint169 = 0;
    end
  end
end


string linebuf170 = "";
logic hitMadPrint170 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc170_inst_done && ((spc170_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint170 = 1;
       linebuf170 = {linebuf170, spc170_phy_pc_w[8:1]};
       if (spc170_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 170, linebuf170);
          linebuf170 = "";
       end
    end else begin
       hitMadPrint170 = 0;
    end
  end
end


string linebuf171 = "";
logic hitMadPrint171 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc171_inst_done && ((spc171_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint171 = 1;
       linebuf171 = {linebuf171, spc171_phy_pc_w[8:1]};
       if (spc171_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 171, linebuf171);
          linebuf171 = "";
       end
    end else begin
       hitMadPrint171 = 0;
    end
  end
end


string linebuf172 = "";
logic hitMadPrint172 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc172_inst_done && ((spc172_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint172 = 1;
       linebuf172 = {linebuf172, spc172_phy_pc_w[8:1]};
       if (spc172_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 172, linebuf172);
          linebuf172 = "";
       end
    end else begin
       hitMadPrint172 = 0;
    end
  end
end


string linebuf173 = "";
logic hitMadPrint173 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc173_inst_done && ((spc173_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint173 = 1;
       linebuf173 = {linebuf173, spc173_phy_pc_w[8:1]};
       if (spc173_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 173, linebuf173);
          linebuf173 = "";
       end
    end else begin
       hitMadPrint173 = 0;
    end
  end
end


string linebuf174 = "";
logic hitMadPrint174 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc174_inst_done && ((spc174_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint174 = 1;
       linebuf174 = {linebuf174, spc174_phy_pc_w[8:1]};
       if (spc174_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 174, linebuf174);
          linebuf174 = "";
       end
    end else begin
       hitMadPrint174 = 0;
    end
  end
end


string linebuf175 = "";
logic hitMadPrint175 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc175_inst_done && ((spc175_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint175 = 1;
       linebuf175 = {linebuf175, spc175_phy_pc_w[8:1]};
       if (spc175_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 175, linebuf175);
          linebuf175 = "";
       end
    end else begin
       hitMadPrint175 = 0;
    end
  end
end


string linebuf176 = "";
logic hitMadPrint176 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc176_inst_done && ((spc176_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint176 = 1;
       linebuf176 = {linebuf176, spc176_phy_pc_w[8:1]};
       if (spc176_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 176, linebuf176);
          linebuf176 = "";
       end
    end else begin
       hitMadPrint176 = 0;
    end
  end
end


string linebuf177 = "";
logic hitMadPrint177 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc177_inst_done && ((spc177_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint177 = 1;
       linebuf177 = {linebuf177, spc177_phy_pc_w[8:1]};
       if (spc177_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 177, linebuf177);
          linebuf177 = "";
       end
    end else begin
       hitMadPrint177 = 0;
    end
  end
end


string linebuf178 = "";
logic hitMadPrint178 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc178_inst_done && ((spc178_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint178 = 1;
       linebuf178 = {linebuf178, spc178_phy_pc_w[8:1]};
       if (spc178_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 178, linebuf178);
          linebuf178 = "";
       end
    end else begin
       hitMadPrint178 = 0;
    end
  end
end


string linebuf179 = "";
logic hitMadPrint179 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc179_inst_done && ((spc179_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint179 = 1;
       linebuf179 = {linebuf179, spc179_phy_pc_w[8:1]};
       if (spc179_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 179, linebuf179);
          linebuf179 = "";
       end
    end else begin
       hitMadPrint179 = 0;
    end
  end
end


string linebuf180 = "";
logic hitMadPrint180 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc180_inst_done && ((spc180_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint180 = 1;
       linebuf180 = {linebuf180, spc180_phy_pc_w[8:1]};
       if (spc180_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 180, linebuf180);
          linebuf180 = "";
       end
    end else begin
       hitMadPrint180 = 0;
    end
  end
end


string linebuf181 = "";
logic hitMadPrint181 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc181_inst_done && ((spc181_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint181 = 1;
       linebuf181 = {linebuf181, spc181_phy_pc_w[8:1]};
       if (spc181_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 181, linebuf181);
          linebuf181 = "";
       end
    end else begin
       hitMadPrint181 = 0;
    end
  end
end


string linebuf182 = "";
logic hitMadPrint182 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc182_inst_done && ((spc182_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint182 = 1;
       linebuf182 = {linebuf182, spc182_phy_pc_w[8:1]};
       if (spc182_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 182, linebuf182);
          linebuf182 = "";
       end
    end else begin
       hitMadPrint182 = 0;
    end
  end
end


string linebuf183 = "";
logic hitMadPrint183 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc183_inst_done && ((spc183_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint183 = 1;
       linebuf183 = {linebuf183, spc183_phy_pc_w[8:1]};
       if (spc183_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 183, linebuf183);
          linebuf183 = "";
       end
    end else begin
       hitMadPrint183 = 0;
    end
  end
end


string linebuf184 = "";
logic hitMadPrint184 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc184_inst_done && ((spc184_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint184 = 1;
       linebuf184 = {linebuf184, spc184_phy_pc_w[8:1]};
       if (spc184_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 184, linebuf184);
          linebuf184 = "";
       end
    end else begin
       hitMadPrint184 = 0;
    end
  end
end


string linebuf185 = "";
logic hitMadPrint185 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc185_inst_done && ((spc185_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint185 = 1;
       linebuf185 = {linebuf185, spc185_phy_pc_w[8:1]};
       if (spc185_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 185, linebuf185);
          linebuf185 = "";
       end
    end else begin
       hitMadPrint185 = 0;
    end
  end
end


string linebuf186 = "";
logic hitMadPrint186 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc186_inst_done && ((spc186_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint186 = 1;
       linebuf186 = {linebuf186, spc186_phy_pc_w[8:1]};
       if (spc186_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 186, linebuf186);
          linebuf186 = "";
       end
    end else begin
       hitMadPrint186 = 0;
    end
  end
end


string linebuf187 = "";
logic hitMadPrint187 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc187_inst_done && ((spc187_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint187 = 1;
       linebuf187 = {linebuf187, spc187_phy_pc_w[8:1]};
       if (spc187_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 187, linebuf187);
          linebuf187 = "";
       end
    end else begin
       hitMadPrint187 = 0;
    end
  end
end


string linebuf188 = "";
logic hitMadPrint188 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc188_inst_done && ((spc188_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint188 = 1;
       linebuf188 = {linebuf188, spc188_phy_pc_w[8:1]};
       if (spc188_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 188, linebuf188);
          linebuf188 = "";
       end
    end else begin
       hitMadPrint188 = 0;
    end
  end
end


string linebuf189 = "";
logic hitMadPrint189 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc189_inst_done && ((spc189_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint189 = 1;
       linebuf189 = {linebuf189, spc189_phy_pc_w[8:1]};
       if (spc189_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 189, linebuf189);
          linebuf189 = "";
       end
    end else begin
       hitMadPrint189 = 0;
    end
  end
end


string linebuf190 = "";
logic hitMadPrint190 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc190_inst_done && ((spc190_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint190 = 1;
       linebuf190 = {linebuf190, spc190_phy_pc_w[8:1]};
       if (spc190_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 190, linebuf190);
          linebuf190 = "";
       end
    end else begin
       hitMadPrint190 = 0;
    end
  end
end


string linebuf191 = "";
logic hitMadPrint191 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc191_inst_done && ((spc191_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint191 = 1;
       linebuf191 = {linebuf191, spc191_phy_pc_w[8:1]};
       if (spc191_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 191, linebuf191);
          linebuf191 = "";
       end
    end else begin
       hitMadPrint191 = 0;
    end
  end
end


string linebuf192 = "";
logic hitMadPrint192 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc192_inst_done && ((spc192_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint192 = 1;
       linebuf192 = {linebuf192, spc192_phy_pc_w[8:1]};
       if (spc192_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 192, linebuf192);
          linebuf192 = "";
       end
    end else begin
       hitMadPrint192 = 0;
    end
  end
end


string linebuf193 = "";
logic hitMadPrint193 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc193_inst_done && ((spc193_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint193 = 1;
       linebuf193 = {linebuf193, spc193_phy_pc_w[8:1]};
       if (spc193_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 193, linebuf193);
          linebuf193 = "";
       end
    end else begin
       hitMadPrint193 = 0;
    end
  end
end


string linebuf194 = "";
logic hitMadPrint194 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc194_inst_done && ((spc194_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint194 = 1;
       linebuf194 = {linebuf194, spc194_phy_pc_w[8:1]};
       if (spc194_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 194, linebuf194);
          linebuf194 = "";
       end
    end else begin
       hitMadPrint194 = 0;
    end
  end
end


string linebuf195 = "";
logic hitMadPrint195 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc195_inst_done && ((spc195_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint195 = 1;
       linebuf195 = {linebuf195, spc195_phy_pc_w[8:1]};
       if (spc195_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 195, linebuf195);
          linebuf195 = "";
       end
    end else begin
       hitMadPrint195 = 0;
    end
  end
end


string linebuf196 = "";
logic hitMadPrint196 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc196_inst_done && ((spc196_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint196 = 1;
       linebuf196 = {linebuf196, spc196_phy_pc_w[8:1]};
       if (spc196_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 196, linebuf196);
          linebuf196 = "";
       end
    end else begin
       hitMadPrint196 = 0;
    end
  end
end


string linebuf197 = "";
logic hitMadPrint197 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc197_inst_done && ((spc197_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint197 = 1;
       linebuf197 = {linebuf197, spc197_phy_pc_w[8:1]};
       if (spc197_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 197, linebuf197);
          linebuf197 = "";
       end
    end else begin
       hitMadPrint197 = 0;
    end
  end
end


string linebuf198 = "";
logic hitMadPrint198 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc198_inst_done && ((spc198_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint198 = 1;
       linebuf198 = {linebuf198, spc198_phy_pc_w[8:1]};
       if (spc198_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 198, linebuf198);
          linebuf198 = "";
       end
    end else begin
       hitMadPrint198 = 0;
    end
  end
end


string linebuf199 = "";
logic hitMadPrint199 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc199_inst_done && ((spc199_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint199 = 1;
       linebuf199 = {linebuf199, spc199_phy_pc_w[8:1]};
       if (spc199_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 199, linebuf199);
          linebuf199 = "";
       end
    end else begin
       hitMadPrint199 = 0;
    end
  end
end


string linebuf200 = "";
logic hitMadPrint200 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc200_inst_done && ((spc200_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint200 = 1;
       linebuf200 = {linebuf200, spc200_phy_pc_w[8:1]};
       if (spc200_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 200, linebuf200);
          linebuf200 = "";
       end
    end else begin
       hitMadPrint200 = 0;
    end
  end
end


string linebuf201 = "";
logic hitMadPrint201 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc201_inst_done && ((spc201_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint201 = 1;
       linebuf201 = {linebuf201, spc201_phy_pc_w[8:1]};
       if (spc201_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 201, linebuf201);
          linebuf201 = "";
       end
    end else begin
       hitMadPrint201 = 0;
    end
  end
end


string linebuf202 = "";
logic hitMadPrint202 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc202_inst_done && ((spc202_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint202 = 1;
       linebuf202 = {linebuf202, spc202_phy_pc_w[8:1]};
       if (spc202_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 202, linebuf202);
          linebuf202 = "";
       end
    end else begin
       hitMadPrint202 = 0;
    end
  end
end


string linebuf203 = "";
logic hitMadPrint203 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc203_inst_done && ((spc203_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint203 = 1;
       linebuf203 = {linebuf203, spc203_phy_pc_w[8:1]};
       if (spc203_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 203, linebuf203);
          linebuf203 = "";
       end
    end else begin
       hitMadPrint203 = 0;
    end
  end
end


string linebuf204 = "";
logic hitMadPrint204 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc204_inst_done && ((spc204_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint204 = 1;
       linebuf204 = {linebuf204, spc204_phy_pc_w[8:1]};
       if (spc204_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 204, linebuf204);
          linebuf204 = "";
       end
    end else begin
       hitMadPrint204 = 0;
    end
  end
end


string linebuf205 = "";
logic hitMadPrint205 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc205_inst_done && ((spc205_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint205 = 1;
       linebuf205 = {linebuf205, spc205_phy_pc_w[8:1]};
       if (spc205_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 205, linebuf205);
          linebuf205 = "";
       end
    end else begin
       hitMadPrint205 = 0;
    end
  end
end


string linebuf206 = "";
logic hitMadPrint206 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc206_inst_done && ((spc206_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint206 = 1;
       linebuf206 = {linebuf206, spc206_phy_pc_w[8:1]};
       if (spc206_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 206, linebuf206);
          linebuf206 = "";
       end
    end else begin
       hitMadPrint206 = 0;
    end
  end
end


string linebuf207 = "";
logic hitMadPrint207 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc207_inst_done && ((spc207_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint207 = 1;
       linebuf207 = {linebuf207, spc207_phy_pc_w[8:1]};
       if (spc207_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 207, linebuf207);
          linebuf207 = "";
       end
    end else begin
       hitMadPrint207 = 0;
    end
  end
end


string linebuf208 = "";
logic hitMadPrint208 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc208_inst_done && ((spc208_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint208 = 1;
       linebuf208 = {linebuf208, spc208_phy_pc_w[8:1]};
       if (spc208_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 208, linebuf208);
          linebuf208 = "";
       end
    end else begin
       hitMadPrint208 = 0;
    end
  end
end


string linebuf209 = "";
logic hitMadPrint209 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc209_inst_done && ((spc209_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint209 = 1;
       linebuf209 = {linebuf209, spc209_phy_pc_w[8:1]};
       if (spc209_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 209, linebuf209);
          linebuf209 = "";
       end
    end else begin
       hitMadPrint209 = 0;
    end
  end
end


string linebuf210 = "";
logic hitMadPrint210 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc210_inst_done && ((spc210_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint210 = 1;
       linebuf210 = {linebuf210, spc210_phy_pc_w[8:1]};
       if (spc210_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 210, linebuf210);
          linebuf210 = "";
       end
    end else begin
       hitMadPrint210 = 0;
    end
  end
end


string linebuf211 = "";
logic hitMadPrint211 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc211_inst_done && ((spc211_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint211 = 1;
       linebuf211 = {linebuf211, spc211_phy_pc_w[8:1]};
       if (spc211_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 211, linebuf211);
          linebuf211 = "";
       end
    end else begin
       hitMadPrint211 = 0;
    end
  end
end


string linebuf212 = "";
logic hitMadPrint212 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc212_inst_done && ((spc212_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint212 = 1;
       linebuf212 = {linebuf212, spc212_phy_pc_w[8:1]};
       if (spc212_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 212, linebuf212);
          linebuf212 = "";
       end
    end else begin
       hitMadPrint212 = 0;
    end
  end
end


string linebuf213 = "";
logic hitMadPrint213 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc213_inst_done && ((spc213_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint213 = 1;
       linebuf213 = {linebuf213, spc213_phy_pc_w[8:1]};
       if (spc213_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 213, linebuf213);
          linebuf213 = "";
       end
    end else begin
       hitMadPrint213 = 0;
    end
  end
end


string linebuf214 = "";
logic hitMadPrint214 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc214_inst_done && ((spc214_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint214 = 1;
       linebuf214 = {linebuf214, spc214_phy_pc_w[8:1]};
       if (spc214_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 214, linebuf214);
          linebuf214 = "";
       end
    end else begin
       hitMadPrint214 = 0;
    end
  end
end


string linebuf215 = "";
logic hitMadPrint215 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc215_inst_done && ((spc215_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint215 = 1;
       linebuf215 = {linebuf215, spc215_phy_pc_w[8:1]};
       if (spc215_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 215, linebuf215);
          linebuf215 = "";
       end
    end else begin
       hitMadPrint215 = 0;
    end
  end
end


string linebuf216 = "";
logic hitMadPrint216 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc216_inst_done && ((spc216_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint216 = 1;
       linebuf216 = {linebuf216, spc216_phy_pc_w[8:1]};
       if (spc216_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 216, linebuf216);
          linebuf216 = "";
       end
    end else begin
       hitMadPrint216 = 0;
    end
  end
end


string linebuf217 = "";
logic hitMadPrint217 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc217_inst_done && ((spc217_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint217 = 1;
       linebuf217 = {linebuf217, spc217_phy_pc_w[8:1]};
       if (spc217_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 217, linebuf217);
          linebuf217 = "";
       end
    end else begin
       hitMadPrint217 = 0;
    end
  end
end


string linebuf218 = "";
logic hitMadPrint218 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc218_inst_done && ((spc218_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint218 = 1;
       linebuf218 = {linebuf218, spc218_phy_pc_w[8:1]};
       if (spc218_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 218, linebuf218);
          linebuf218 = "";
       end
    end else begin
       hitMadPrint218 = 0;
    end
  end
end


string linebuf219 = "";
logic hitMadPrint219 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc219_inst_done && ((spc219_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint219 = 1;
       linebuf219 = {linebuf219, spc219_phy_pc_w[8:1]};
       if (spc219_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 219, linebuf219);
          linebuf219 = "";
       end
    end else begin
       hitMadPrint219 = 0;
    end
  end
end


string linebuf220 = "";
logic hitMadPrint220 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc220_inst_done && ((spc220_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint220 = 1;
       linebuf220 = {linebuf220, spc220_phy_pc_w[8:1]};
       if (spc220_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 220, linebuf220);
          linebuf220 = "";
       end
    end else begin
       hitMadPrint220 = 0;
    end
  end
end


string linebuf221 = "";
logic hitMadPrint221 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc221_inst_done && ((spc221_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint221 = 1;
       linebuf221 = {linebuf221, spc221_phy_pc_w[8:1]};
       if (spc221_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 221, linebuf221);
          linebuf221 = "";
       end
    end else begin
       hitMadPrint221 = 0;
    end
  end
end


string linebuf222 = "";
logic hitMadPrint222 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc222_inst_done && ((spc222_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint222 = 1;
       linebuf222 = {linebuf222, spc222_phy_pc_w[8:1]};
       if (spc222_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 222, linebuf222);
          linebuf222 = "";
       end
    end else begin
       hitMadPrint222 = 0;
    end
  end
end


string linebuf223 = "";
logic hitMadPrint223 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc223_inst_done && ((spc223_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint223 = 1;
       linebuf223 = {linebuf223, spc223_phy_pc_w[8:1]};
       if (spc223_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 223, linebuf223);
          linebuf223 = "";
       end
    end else begin
       hitMadPrint223 = 0;
    end
  end
end


string linebuf224 = "";
logic hitMadPrint224 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc224_inst_done && ((spc224_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint224 = 1;
       linebuf224 = {linebuf224, spc224_phy_pc_w[8:1]};
       if (spc224_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 224, linebuf224);
          linebuf224 = "";
       end
    end else begin
       hitMadPrint224 = 0;
    end
  end
end


string linebuf225 = "";
logic hitMadPrint225 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc225_inst_done && ((spc225_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint225 = 1;
       linebuf225 = {linebuf225, spc225_phy_pc_w[8:1]};
       if (spc225_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 225, linebuf225);
          linebuf225 = "";
       end
    end else begin
       hitMadPrint225 = 0;
    end
  end
end


string linebuf226 = "";
logic hitMadPrint226 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc226_inst_done && ((spc226_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint226 = 1;
       linebuf226 = {linebuf226, spc226_phy_pc_w[8:1]};
       if (spc226_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 226, linebuf226);
          linebuf226 = "";
       end
    end else begin
       hitMadPrint226 = 0;
    end
  end
end


string linebuf227 = "";
logic hitMadPrint227 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc227_inst_done && ((spc227_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint227 = 1;
       linebuf227 = {linebuf227, spc227_phy_pc_w[8:1]};
       if (spc227_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 227, linebuf227);
          linebuf227 = "";
       end
    end else begin
       hitMadPrint227 = 0;
    end
  end
end


string linebuf228 = "";
logic hitMadPrint228 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc228_inst_done && ((spc228_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint228 = 1;
       linebuf228 = {linebuf228, spc228_phy_pc_w[8:1]};
       if (spc228_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 228, linebuf228);
          linebuf228 = "";
       end
    end else begin
       hitMadPrint228 = 0;
    end
  end
end


string linebuf229 = "";
logic hitMadPrint229 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc229_inst_done && ((spc229_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint229 = 1;
       linebuf229 = {linebuf229, spc229_phy_pc_w[8:1]};
       if (spc229_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 229, linebuf229);
          linebuf229 = "";
       end
    end else begin
       hitMadPrint229 = 0;
    end
  end
end


string linebuf230 = "";
logic hitMadPrint230 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc230_inst_done && ((spc230_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint230 = 1;
       linebuf230 = {linebuf230, spc230_phy_pc_w[8:1]};
       if (spc230_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 230, linebuf230);
          linebuf230 = "";
       end
    end else begin
       hitMadPrint230 = 0;
    end
  end
end


string linebuf231 = "";
logic hitMadPrint231 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc231_inst_done && ((spc231_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint231 = 1;
       linebuf231 = {linebuf231, spc231_phy_pc_w[8:1]};
       if (spc231_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 231, linebuf231);
          linebuf231 = "";
       end
    end else begin
       hitMadPrint231 = 0;
    end
  end
end


string linebuf232 = "";
logic hitMadPrint232 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc232_inst_done && ((spc232_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint232 = 1;
       linebuf232 = {linebuf232, spc232_phy_pc_w[8:1]};
       if (spc232_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 232, linebuf232);
          linebuf232 = "";
       end
    end else begin
       hitMadPrint232 = 0;
    end
  end
end


string linebuf233 = "";
logic hitMadPrint233 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc233_inst_done && ((spc233_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint233 = 1;
       linebuf233 = {linebuf233, spc233_phy_pc_w[8:1]};
       if (spc233_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 233, linebuf233);
          linebuf233 = "";
       end
    end else begin
       hitMadPrint233 = 0;
    end
  end
end


string linebuf234 = "";
logic hitMadPrint234 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc234_inst_done && ((spc234_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint234 = 1;
       linebuf234 = {linebuf234, spc234_phy_pc_w[8:1]};
       if (spc234_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 234, linebuf234);
          linebuf234 = "";
       end
    end else begin
       hitMadPrint234 = 0;
    end
  end
end


string linebuf235 = "";
logic hitMadPrint235 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc235_inst_done && ((spc235_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint235 = 1;
       linebuf235 = {linebuf235, spc235_phy_pc_w[8:1]};
       if (spc235_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 235, linebuf235);
          linebuf235 = "";
       end
    end else begin
       hitMadPrint235 = 0;
    end
  end
end


string linebuf236 = "";
logic hitMadPrint236 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc236_inst_done && ((spc236_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint236 = 1;
       linebuf236 = {linebuf236, spc236_phy_pc_w[8:1]};
       if (spc236_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 236, linebuf236);
          linebuf236 = "";
       end
    end else begin
       hitMadPrint236 = 0;
    end
  end
end


string linebuf237 = "";
logic hitMadPrint237 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc237_inst_done && ((spc237_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint237 = 1;
       linebuf237 = {linebuf237, spc237_phy_pc_w[8:1]};
       if (spc237_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 237, linebuf237);
          linebuf237 = "";
       end
    end else begin
       hitMadPrint237 = 0;
    end
  end
end


string linebuf238 = "";
logic hitMadPrint238 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc238_inst_done && ((spc238_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint238 = 1;
       linebuf238 = {linebuf238, spc238_phy_pc_w[8:1]};
       if (spc238_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 238, linebuf238);
          linebuf238 = "";
       end
    end else begin
       hitMadPrint238 = 0;
    end
  end
end


string linebuf239 = "";
logic hitMadPrint239 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc239_inst_done && ((spc239_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint239 = 1;
       linebuf239 = {linebuf239, spc239_phy_pc_w[8:1]};
       if (spc239_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 239, linebuf239);
          linebuf239 = "";
       end
    end else begin
       hitMadPrint239 = 0;
    end
  end
end


string linebuf240 = "";
logic hitMadPrint240 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc240_inst_done && ((spc240_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint240 = 1;
       linebuf240 = {linebuf240, spc240_phy_pc_w[8:1]};
       if (spc240_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 240, linebuf240);
          linebuf240 = "";
       end
    end else begin
       hitMadPrint240 = 0;
    end
  end
end


string linebuf241 = "";
logic hitMadPrint241 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc241_inst_done && ((spc241_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint241 = 1;
       linebuf241 = {linebuf241, spc241_phy_pc_w[8:1]};
       if (spc241_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 241, linebuf241);
          linebuf241 = "";
       end
    end else begin
       hitMadPrint241 = 0;
    end
  end
end


string linebuf242 = "";
logic hitMadPrint242 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc242_inst_done && ((spc242_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint242 = 1;
       linebuf242 = {linebuf242, spc242_phy_pc_w[8:1]};
       if (spc242_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 242, linebuf242);
          linebuf242 = "";
       end
    end else begin
       hitMadPrint242 = 0;
    end
  end
end


string linebuf243 = "";
logic hitMadPrint243 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc243_inst_done && ((spc243_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint243 = 1;
       linebuf243 = {linebuf243, spc243_phy_pc_w[8:1]};
       if (spc243_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 243, linebuf243);
          linebuf243 = "";
       end
    end else begin
       hitMadPrint243 = 0;
    end
  end
end


string linebuf244 = "";
logic hitMadPrint244 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc244_inst_done && ((spc244_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint244 = 1;
       linebuf244 = {linebuf244, spc244_phy_pc_w[8:1]};
       if (spc244_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 244, linebuf244);
          linebuf244 = "";
       end
    end else begin
       hitMadPrint244 = 0;
    end
  end
end


string linebuf245 = "";
logic hitMadPrint245 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc245_inst_done && ((spc245_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint245 = 1;
       linebuf245 = {linebuf245, spc245_phy_pc_w[8:1]};
       if (spc245_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 245, linebuf245);
          linebuf245 = "";
       end
    end else begin
       hitMadPrint245 = 0;
    end
  end
end


string linebuf246 = "";
logic hitMadPrint246 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc246_inst_done && ((spc246_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint246 = 1;
       linebuf246 = {linebuf246, spc246_phy_pc_w[8:1]};
       if (spc246_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 246, linebuf246);
          linebuf246 = "";
       end
    end else begin
       hitMadPrint246 = 0;
    end
  end
end


string linebuf247 = "";
logic hitMadPrint247 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc247_inst_done && ((spc247_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint247 = 1;
       linebuf247 = {linebuf247, spc247_phy_pc_w[8:1]};
       if (spc247_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 247, linebuf247);
          linebuf247 = "";
       end
    end else begin
       hitMadPrint247 = 0;
    end
  end
end


string linebuf248 = "";
logic hitMadPrint248 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc248_inst_done && ((spc248_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint248 = 1;
       linebuf248 = {linebuf248, spc248_phy_pc_w[8:1]};
       if (spc248_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 248, linebuf248);
          linebuf248 = "";
       end
    end else begin
       hitMadPrint248 = 0;
    end
  end
end


string linebuf249 = "";
logic hitMadPrint249 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc249_inst_done && ((spc249_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint249 = 1;
       linebuf249 = {linebuf249, spc249_phy_pc_w[8:1]};
       if (spc249_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 249, linebuf249);
          linebuf249 = "";
       end
    end else begin
       hitMadPrint249 = 0;
    end
  end
end


string linebuf250 = "";
logic hitMadPrint250 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc250_inst_done && ((spc250_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint250 = 1;
       linebuf250 = {linebuf250, spc250_phy_pc_w[8:1]};
       if (spc250_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 250, linebuf250);
          linebuf250 = "";
       end
    end else begin
       hitMadPrint250 = 0;
    end
  end
end


string linebuf251 = "";
logic hitMadPrint251 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc251_inst_done && ((spc251_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint251 = 1;
       linebuf251 = {linebuf251, spc251_phy_pc_w[8:1]};
       if (spc251_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 251, linebuf251);
          linebuf251 = "";
       end
    end else begin
       hitMadPrint251 = 0;
    end
  end
end


string linebuf252 = "";
logic hitMadPrint252 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc252_inst_done && ((spc252_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint252 = 1;
       linebuf252 = {linebuf252, spc252_phy_pc_w[8:1]};
       if (spc252_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 252, linebuf252);
          linebuf252 = "";
       end
    end else begin
       hitMadPrint252 = 0;
    end
  end
end


string linebuf253 = "";
logic hitMadPrint253 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc253_inst_done && ((spc253_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint253 = 1;
       linebuf253 = {linebuf253, spc253_phy_pc_w[8:1]};
       if (spc253_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 253, linebuf253);
          linebuf253 = "";
       end
    end else begin
       hitMadPrint253 = 0;
    end
  end
end


string linebuf254 = "";
logic hitMadPrint254 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc254_inst_done && ((spc254_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint254 = 1;
       linebuf254 = {linebuf254, spc254_phy_pc_w[8:1]};
       if (spc254_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 254, linebuf254);
          linebuf254 = "";
       end
    end else begin
       hitMadPrint254 = 0;
    end
  end
end


string linebuf255 = "";
logic hitMadPrint255 = 0;
always @(posedge clk) begin
  if (rst_l) begin
    if (spc255_inst_done && ((spc255_phy_pc_w >> 9) == (64'h80000400 >> 9))) begin
       hitMadPrint255 = 1;
       linebuf255 = {linebuf255, spc255_phy_pc_w[8:1]};
       if (spc255_phy_pc_w[8:1] == "\n") begin
          $write("%016t hart %4d: %s", $time, 255, linebuf255);
          linebuf255 = "";
       end
    end else begin
       hitMadPrint255 = 0;
    end
  end
end




//main routine of pc cmp to finish the simulation.
always @(posedge clk)begin
    if(rst_l)begin
        if(|done[`PITON_NUM_TILES-1:0]) begin

        if (done[0]) begin
            timeout[long_cpuid0] = 0;
            //check_bad_trap(spc0_phy_pc_w, 0, long_cpuid0);
            if(active_thread[long_cpuid0])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc0_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid0/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 0 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid0]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc0_phy_pc_w))
                begin
                    if(good[long_cpuid0/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid0 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid0/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid0])
        end // if (done[0])

        if (done[1]) begin
            timeout[long_cpuid1] = 0;
            //check_bad_trap(spc1_phy_pc_w, 1, long_cpuid1);
            if(active_thread[long_cpuid1])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc1_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid1/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 1 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid1]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc1_phy_pc_w))
                begin
                    if(good[long_cpuid1/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid1 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid1/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid1])
        end // if (done[1])

        if (done[2]) begin
            timeout[long_cpuid2] = 0;
            //check_bad_trap(spc2_phy_pc_w, 2, long_cpuid2);
            if(active_thread[long_cpuid2])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc2_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid2/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 2 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid2]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc2_phy_pc_w))
                begin
                    if(good[long_cpuid2/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid2 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid2/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid2])
        end // if (done[2])

        if (done[3]) begin
            timeout[long_cpuid3] = 0;
            //check_bad_trap(spc3_phy_pc_w, 3, long_cpuid3);
            if(active_thread[long_cpuid3])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc3_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid3/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 3 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid3]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc3_phy_pc_w))
                begin
                    if(good[long_cpuid3/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid3 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid3/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid3])
        end // if (done[3])

        if (done[4]) begin
            timeout[long_cpuid4] = 0;
            //check_bad_trap(spc4_phy_pc_w, 4, long_cpuid4);
            if(active_thread[long_cpuid4])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc4_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid4/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 4 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid4]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc4_phy_pc_w))
                begin
                    if(good[long_cpuid4/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid4 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid4/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid4])
        end // if (done[4])

        if (done[5]) begin
            timeout[long_cpuid5] = 0;
            //check_bad_trap(spc5_phy_pc_w, 5, long_cpuid5);
            if(active_thread[long_cpuid5])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc5_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid5/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 5 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid5]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc5_phy_pc_w))
                begin
                    if(good[long_cpuid5/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid5 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid5/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid5])
        end // if (done[5])

        if (done[6]) begin
            timeout[long_cpuid6] = 0;
            //check_bad_trap(spc6_phy_pc_w, 6, long_cpuid6);
            if(active_thread[long_cpuid6])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc6_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid6/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 6 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid6]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc6_phy_pc_w))
                begin
                    if(good[long_cpuid6/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid6 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid6/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid6])
        end // if (done[6])

        if (done[7]) begin
            timeout[long_cpuid7] = 0;
            //check_bad_trap(spc7_phy_pc_w, 7, long_cpuid7);
            if(active_thread[long_cpuid7])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc7_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid7/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 7 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid7]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc7_phy_pc_w))
                begin
                    if(good[long_cpuid7/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid7 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid7/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid7])
        end // if (done[7])

        if (done[8]) begin
            timeout[long_cpuid8] = 0;
            //check_bad_trap(spc8_phy_pc_w, 8, long_cpuid8);
            if(active_thread[long_cpuid8])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc8_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid8/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 8 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid8]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc8_phy_pc_w))
                begin
                    if(good[long_cpuid8/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid8 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid8/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid8])
        end // if (done[8])

        if (done[9]) begin
            timeout[long_cpuid9] = 0;
            //check_bad_trap(spc9_phy_pc_w, 9, long_cpuid9);
            if(active_thread[long_cpuid9])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc9_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid9/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 9 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid9]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc9_phy_pc_w))
                begin
                    if(good[long_cpuid9/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid9 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid9/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid9])
        end // if (done[9])

        if (done[10]) begin
            timeout[long_cpuid10] = 0;
            //check_bad_trap(spc10_phy_pc_w, 10, long_cpuid10);
            if(active_thread[long_cpuid10])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc10_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid10/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 10 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid10]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc10_phy_pc_w))
                begin
                    if(good[long_cpuid10/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid10 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid10/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid10])
        end // if (done[10])

        if (done[11]) begin
            timeout[long_cpuid11] = 0;
            //check_bad_trap(spc11_phy_pc_w, 11, long_cpuid11);
            if(active_thread[long_cpuid11])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc11_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid11/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 11 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid11]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc11_phy_pc_w))
                begin
                    if(good[long_cpuid11/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid11 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid11/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid11])
        end // if (done[11])

        if (done[12]) begin
            timeout[long_cpuid12] = 0;
            //check_bad_trap(spc12_phy_pc_w, 12, long_cpuid12);
            if(active_thread[long_cpuid12])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc12_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid12/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 12 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid12]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc12_phy_pc_w))
                begin
                    if(good[long_cpuid12/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid12 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid12/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid12])
        end // if (done[12])

        if (done[13]) begin
            timeout[long_cpuid13] = 0;
            //check_bad_trap(spc13_phy_pc_w, 13, long_cpuid13);
            if(active_thread[long_cpuid13])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc13_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid13/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 13 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid13]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc13_phy_pc_w))
                begin
                    if(good[long_cpuid13/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid13 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid13/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid13])
        end // if (done[13])

        if (done[14]) begin
            timeout[long_cpuid14] = 0;
            //check_bad_trap(spc14_phy_pc_w, 14, long_cpuid14);
            if(active_thread[long_cpuid14])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc14_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid14/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 14 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid14]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc14_phy_pc_w))
                begin
                    if(good[long_cpuid14/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid14 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid14/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid14])
        end // if (done[14])

        if (done[15]) begin
            timeout[long_cpuid15] = 0;
            //check_bad_trap(spc15_phy_pc_w, 15, long_cpuid15);
            if(active_thread[long_cpuid15])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc15_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid15/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 15 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid15]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc15_phy_pc_w))
                begin
                    if(good[long_cpuid15/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid15 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid15/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid15])
        end // if (done[15])

        if (done[16]) begin
            timeout[long_cpuid16] = 0;
            //check_bad_trap(spc16_phy_pc_w, 16, long_cpuid16);
            if(active_thread[long_cpuid16])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc16_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid16/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 16 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid16]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc16_phy_pc_w))
                begin
                    if(good[long_cpuid16/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid16 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid16/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid16])
        end // if (done[16])

        if (done[17]) begin
            timeout[long_cpuid17] = 0;
            //check_bad_trap(spc17_phy_pc_w, 17, long_cpuid17);
            if(active_thread[long_cpuid17])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc17_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid17/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 17 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid17]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc17_phy_pc_w))
                begin
                    if(good[long_cpuid17/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid17 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid17/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid17])
        end // if (done[17])

        if (done[18]) begin
            timeout[long_cpuid18] = 0;
            //check_bad_trap(spc18_phy_pc_w, 18, long_cpuid18);
            if(active_thread[long_cpuid18])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc18_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid18/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 18 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid18]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc18_phy_pc_w))
                begin
                    if(good[long_cpuid18/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid18 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid18/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid18])
        end // if (done[18])

        if (done[19]) begin
            timeout[long_cpuid19] = 0;
            //check_bad_trap(spc19_phy_pc_w, 19, long_cpuid19);
            if(active_thread[long_cpuid19])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc19_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid19/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 19 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid19]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc19_phy_pc_w))
                begin
                    if(good[long_cpuid19/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid19 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid19/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid19])
        end // if (done[19])

        if (done[20]) begin
            timeout[long_cpuid20] = 0;
            //check_bad_trap(spc20_phy_pc_w, 20, long_cpuid20);
            if(active_thread[long_cpuid20])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc20_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid20/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 20 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid20]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc20_phy_pc_w))
                begin
                    if(good[long_cpuid20/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid20 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid20/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid20])
        end // if (done[20])

        if (done[21]) begin
            timeout[long_cpuid21] = 0;
            //check_bad_trap(spc21_phy_pc_w, 21, long_cpuid21);
            if(active_thread[long_cpuid21])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc21_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid21/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 21 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid21]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc21_phy_pc_w))
                begin
                    if(good[long_cpuid21/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid21 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid21/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid21])
        end // if (done[21])

        if (done[22]) begin
            timeout[long_cpuid22] = 0;
            //check_bad_trap(spc22_phy_pc_w, 22, long_cpuid22);
            if(active_thread[long_cpuid22])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc22_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid22/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 22 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid22]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc22_phy_pc_w))
                begin
                    if(good[long_cpuid22/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid22 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid22/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid22])
        end // if (done[22])

        if (done[23]) begin
            timeout[long_cpuid23] = 0;
            //check_bad_trap(spc23_phy_pc_w, 23, long_cpuid23);
            if(active_thread[long_cpuid23])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc23_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid23/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 23 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid23]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc23_phy_pc_w))
                begin
                    if(good[long_cpuid23/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid23 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid23/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid23])
        end // if (done[23])

        if (done[24]) begin
            timeout[long_cpuid24] = 0;
            //check_bad_trap(spc24_phy_pc_w, 24, long_cpuid24);
            if(active_thread[long_cpuid24])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc24_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid24/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 24 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid24]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc24_phy_pc_w))
                begin
                    if(good[long_cpuid24/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid24 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid24/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid24])
        end // if (done[24])

        if (done[25]) begin
            timeout[long_cpuid25] = 0;
            //check_bad_trap(spc25_phy_pc_w, 25, long_cpuid25);
            if(active_thread[long_cpuid25])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc25_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid25/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 25 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid25]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc25_phy_pc_w))
                begin
                    if(good[long_cpuid25/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid25 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid25/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid25])
        end // if (done[25])

        if (done[26]) begin
            timeout[long_cpuid26] = 0;
            //check_bad_trap(spc26_phy_pc_w, 26, long_cpuid26);
            if(active_thread[long_cpuid26])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc26_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid26/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 26 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid26]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc26_phy_pc_w))
                begin
                    if(good[long_cpuid26/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid26 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid26/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid26])
        end // if (done[26])

        if (done[27]) begin
            timeout[long_cpuid27] = 0;
            //check_bad_trap(spc27_phy_pc_w, 27, long_cpuid27);
            if(active_thread[long_cpuid27])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc27_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid27/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 27 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid27]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc27_phy_pc_w))
                begin
                    if(good[long_cpuid27/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid27 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid27/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid27])
        end // if (done[27])

        if (done[28]) begin
            timeout[long_cpuid28] = 0;
            //check_bad_trap(spc28_phy_pc_w, 28, long_cpuid28);
            if(active_thread[long_cpuid28])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc28_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid28/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 28 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid28]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc28_phy_pc_w))
                begin
                    if(good[long_cpuid28/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid28 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid28/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid28])
        end // if (done[28])

        if (done[29]) begin
            timeout[long_cpuid29] = 0;
            //check_bad_trap(spc29_phy_pc_w, 29, long_cpuid29);
            if(active_thread[long_cpuid29])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc29_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid29/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 29 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid29]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc29_phy_pc_w))
                begin
                    if(good[long_cpuid29/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid29 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid29/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid29])
        end // if (done[29])

        if (done[30]) begin
            timeout[long_cpuid30] = 0;
            //check_bad_trap(spc30_phy_pc_w, 30, long_cpuid30);
            if(active_thread[long_cpuid30])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc30_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid30/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 30 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid30]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc30_phy_pc_w))
                begin
                    if(good[long_cpuid30/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid30 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid30/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid30])
        end // if (done[30])

        if (done[31]) begin
            timeout[long_cpuid31] = 0;
            //check_bad_trap(spc31_phy_pc_w, 31, long_cpuid31);
            if(active_thread[long_cpuid31])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc31_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid31/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 31 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid31]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc31_phy_pc_w))
                begin
                    if(good[long_cpuid31/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid31 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid31/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid31])
        end // if (done[31])

        if (done[32]) begin
            timeout[long_cpuid32] = 0;
            //check_bad_trap(spc32_phy_pc_w, 32, long_cpuid32);
            if(active_thread[long_cpuid32])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc32_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid32/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 32 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid32]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc32_phy_pc_w))
                begin
                    if(good[long_cpuid32/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid32 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid32/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid32])
        end // if (done[32])

        if (done[33]) begin
            timeout[long_cpuid33] = 0;
            //check_bad_trap(spc33_phy_pc_w, 33, long_cpuid33);
            if(active_thread[long_cpuid33])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc33_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid33/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 33 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid33]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc33_phy_pc_w))
                begin
                    if(good[long_cpuid33/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid33 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid33/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid33])
        end // if (done[33])

        if (done[34]) begin
            timeout[long_cpuid34] = 0;
            //check_bad_trap(spc34_phy_pc_w, 34, long_cpuid34);
            if(active_thread[long_cpuid34])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc34_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid34/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 34 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid34]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc34_phy_pc_w))
                begin
                    if(good[long_cpuid34/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid34 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid34/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid34])
        end // if (done[34])

        if (done[35]) begin
            timeout[long_cpuid35] = 0;
            //check_bad_trap(spc35_phy_pc_w, 35, long_cpuid35);
            if(active_thread[long_cpuid35])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc35_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid35/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 35 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid35]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc35_phy_pc_w))
                begin
                    if(good[long_cpuid35/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid35 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid35/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid35])
        end // if (done[35])

        if (done[36]) begin
            timeout[long_cpuid36] = 0;
            //check_bad_trap(spc36_phy_pc_w, 36, long_cpuid36);
            if(active_thread[long_cpuid36])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc36_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid36/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 36 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid36]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc36_phy_pc_w))
                begin
                    if(good[long_cpuid36/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid36 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid36/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid36])
        end // if (done[36])

        if (done[37]) begin
            timeout[long_cpuid37] = 0;
            //check_bad_trap(spc37_phy_pc_w, 37, long_cpuid37);
            if(active_thread[long_cpuid37])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc37_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid37/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 37 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid37]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc37_phy_pc_w))
                begin
                    if(good[long_cpuid37/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid37 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid37/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid37])
        end // if (done[37])

        if (done[38]) begin
            timeout[long_cpuid38] = 0;
            //check_bad_trap(spc38_phy_pc_w, 38, long_cpuid38);
            if(active_thread[long_cpuid38])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc38_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid38/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 38 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid38]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc38_phy_pc_w))
                begin
                    if(good[long_cpuid38/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid38 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid38/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid38])
        end // if (done[38])

        if (done[39]) begin
            timeout[long_cpuid39] = 0;
            //check_bad_trap(spc39_phy_pc_w, 39, long_cpuid39);
            if(active_thread[long_cpuid39])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc39_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid39/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 39 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid39]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc39_phy_pc_w))
                begin
                    if(good[long_cpuid39/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid39 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid39/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid39])
        end // if (done[39])

        if (done[40]) begin
            timeout[long_cpuid40] = 0;
            //check_bad_trap(spc40_phy_pc_w, 40, long_cpuid40);
            if(active_thread[long_cpuid40])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc40_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid40/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 40 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid40]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc40_phy_pc_w))
                begin
                    if(good[long_cpuid40/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid40 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid40/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid40])
        end // if (done[40])

        if (done[41]) begin
            timeout[long_cpuid41] = 0;
            //check_bad_trap(spc41_phy_pc_w, 41, long_cpuid41);
            if(active_thread[long_cpuid41])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc41_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid41/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 41 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid41]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc41_phy_pc_w))
                begin
                    if(good[long_cpuid41/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid41 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid41/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid41])
        end // if (done[41])

        if (done[42]) begin
            timeout[long_cpuid42] = 0;
            //check_bad_trap(spc42_phy_pc_w, 42, long_cpuid42);
            if(active_thread[long_cpuid42])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc42_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid42/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 42 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid42]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc42_phy_pc_w))
                begin
                    if(good[long_cpuid42/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid42 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid42/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid42])
        end // if (done[42])

        if (done[43]) begin
            timeout[long_cpuid43] = 0;
            //check_bad_trap(spc43_phy_pc_w, 43, long_cpuid43);
            if(active_thread[long_cpuid43])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc43_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid43/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 43 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid43]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc43_phy_pc_w))
                begin
                    if(good[long_cpuid43/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid43 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid43/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid43])
        end // if (done[43])

        if (done[44]) begin
            timeout[long_cpuid44] = 0;
            //check_bad_trap(spc44_phy_pc_w, 44, long_cpuid44);
            if(active_thread[long_cpuid44])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc44_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid44/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 44 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid44]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc44_phy_pc_w))
                begin
                    if(good[long_cpuid44/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid44 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid44/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid44])
        end // if (done[44])

        if (done[45]) begin
            timeout[long_cpuid45] = 0;
            //check_bad_trap(spc45_phy_pc_w, 45, long_cpuid45);
            if(active_thread[long_cpuid45])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc45_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid45/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 45 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid45]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc45_phy_pc_w))
                begin
                    if(good[long_cpuid45/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid45 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid45/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid45])
        end // if (done[45])

        if (done[46]) begin
            timeout[long_cpuid46] = 0;
            //check_bad_trap(spc46_phy_pc_w, 46, long_cpuid46);
            if(active_thread[long_cpuid46])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc46_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid46/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 46 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid46]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc46_phy_pc_w))
                begin
                    if(good[long_cpuid46/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid46 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid46/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid46])
        end // if (done[46])

        if (done[47]) begin
            timeout[long_cpuid47] = 0;
            //check_bad_trap(spc47_phy_pc_w, 47, long_cpuid47);
            if(active_thread[long_cpuid47])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc47_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid47/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 47 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid47]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc47_phy_pc_w))
                begin
                    if(good[long_cpuid47/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid47 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid47/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid47])
        end // if (done[47])

        if (done[48]) begin
            timeout[long_cpuid48] = 0;
            //check_bad_trap(spc48_phy_pc_w, 48, long_cpuid48);
            if(active_thread[long_cpuid48])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc48_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid48/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 48 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid48]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc48_phy_pc_w))
                begin
                    if(good[long_cpuid48/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid48 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid48/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid48])
        end // if (done[48])

        if (done[49]) begin
            timeout[long_cpuid49] = 0;
            //check_bad_trap(spc49_phy_pc_w, 49, long_cpuid49);
            if(active_thread[long_cpuid49])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc49_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid49/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 49 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid49]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc49_phy_pc_w))
                begin
                    if(good[long_cpuid49/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid49 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid49/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid49])
        end // if (done[49])

        if (done[50]) begin
            timeout[long_cpuid50] = 0;
            //check_bad_trap(spc50_phy_pc_w, 50, long_cpuid50);
            if(active_thread[long_cpuid50])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc50_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid50/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 50 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid50]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc50_phy_pc_w))
                begin
                    if(good[long_cpuid50/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid50 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid50/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid50])
        end // if (done[50])

        if (done[51]) begin
            timeout[long_cpuid51] = 0;
            //check_bad_trap(spc51_phy_pc_w, 51, long_cpuid51);
            if(active_thread[long_cpuid51])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc51_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid51/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 51 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid51]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc51_phy_pc_w))
                begin
                    if(good[long_cpuid51/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid51 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid51/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid51])
        end // if (done[51])

        if (done[52]) begin
            timeout[long_cpuid52] = 0;
            //check_bad_trap(spc52_phy_pc_w, 52, long_cpuid52);
            if(active_thread[long_cpuid52])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc52_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid52/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 52 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid52]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc52_phy_pc_w))
                begin
                    if(good[long_cpuid52/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid52 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid52/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid52])
        end // if (done[52])

        if (done[53]) begin
            timeout[long_cpuid53] = 0;
            //check_bad_trap(spc53_phy_pc_w, 53, long_cpuid53);
            if(active_thread[long_cpuid53])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc53_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid53/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 53 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid53]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc53_phy_pc_w))
                begin
                    if(good[long_cpuid53/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid53 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid53/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid53])
        end // if (done[53])

        if (done[54]) begin
            timeout[long_cpuid54] = 0;
            //check_bad_trap(spc54_phy_pc_w, 54, long_cpuid54);
            if(active_thread[long_cpuid54])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc54_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid54/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 54 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid54]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc54_phy_pc_w))
                begin
                    if(good[long_cpuid54/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid54 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid54/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid54])
        end // if (done[54])

        if (done[55]) begin
            timeout[long_cpuid55] = 0;
            //check_bad_trap(spc55_phy_pc_w, 55, long_cpuid55);
            if(active_thread[long_cpuid55])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc55_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid55/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 55 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid55]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc55_phy_pc_w))
                begin
                    if(good[long_cpuid55/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid55 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid55/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid55])
        end // if (done[55])

        if (done[56]) begin
            timeout[long_cpuid56] = 0;
            //check_bad_trap(spc56_phy_pc_w, 56, long_cpuid56);
            if(active_thread[long_cpuid56])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc56_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid56/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 56 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid56]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc56_phy_pc_w))
                begin
                    if(good[long_cpuid56/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid56 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid56/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid56])
        end // if (done[56])

        if (done[57]) begin
            timeout[long_cpuid57] = 0;
            //check_bad_trap(spc57_phy_pc_w, 57, long_cpuid57);
            if(active_thread[long_cpuid57])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc57_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid57/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 57 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid57]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc57_phy_pc_w))
                begin
                    if(good[long_cpuid57/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid57 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid57/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid57])
        end // if (done[57])

        if (done[58]) begin
            timeout[long_cpuid58] = 0;
            //check_bad_trap(spc58_phy_pc_w, 58, long_cpuid58);
            if(active_thread[long_cpuid58])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc58_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid58/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 58 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid58]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc58_phy_pc_w))
                begin
                    if(good[long_cpuid58/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid58 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid58/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid58])
        end // if (done[58])

        if (done[59]) begin
            timeout[long_cpuid59] = 0;
            //check_bad_trap(spc59_phy_pc_w, 59, long_cpuid59);
            if(active_thread[long_cpuid59])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc59_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid59/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 59 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid59]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc59_phy_pc_w))
                begin
                    if(good[long_cpuid59/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid59 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid59/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid59])
        end // if (done[59])

        if (done[60]) begin
            timeout[long_cpuid60] = 0;
            //check_bad_trap(spc60_phy_pc_w, 60, long_cpuid60);
            if(active_thread[long_cpuid60])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc60_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid60/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 60 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid60]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc60_phy_pc_w))
                begin
                    if(good[long_cpuid60/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid60 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid60/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid60])
        end // if (done[60])

        if (done[61]) begin
            timeout[long_cpuid61] = 0;
            //check_bad_trap(spc61_phy_pc_w, 61, long_cpuid61);
            if(active_thread[long_cpuid61])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc61_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid61/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 61 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid61]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc61_phy_pc_w))
                begin
                    if(good[long_cpuid61/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid61 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid61/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid61])
        end // if (done[61])

        if (done[62]) begin
            timeout[long_cpuid62] = 0;
            //check_bad_trap(spc62_phy_pc_w, 62, long_cpuid62);
            if(active_thread[long_cpuid62])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc62_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid62/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 62 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid62]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc62_phy_pc_w))
                begin
                    if(good[long_cpuid62/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid62 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid62/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid62])
        end // if (done[62])

        if (done[63]) begin
            timeout[long_cpuid63] = 0;
            //check_bad_trap(spc63_phy_pc_w, 63, long_cpuid63);
            if(active_thread[long_cpuid63])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc63_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid63/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 63 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid63]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc63_phy_pc_w))
                begin
                    if(good[long_cpuid63/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid63 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid63/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid63])
        end // if (done[63])

        if (done[64]) begin
            timeout[long_cpuid64] = 0;
            //check_bad_trap(spc64_phy_pc_w, 64, long_cpuid64);
            if(active_thread[long_cpuid64])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc64_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid64/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 64 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid64]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc64_phy_pc_w))
                begin
                    if(good[long_cpuid64/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid64 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid64/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid64])
        end // if (done[64])

        if (done[65]) begin
            timeout[long_cpuid65] = 0;
            //check_bad_trap(spc65_phy_pc_w, 65, long_cpuid65);
            if(active_thread[long_cpuid65])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc65_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid65/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 65 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid65]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc65_phy_pc_w))
                begin
                    if(good[long_cpuid65/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid65 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid65/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid65])
        end // if (done[65])

        if (done[66]) begin
            timeout[long_cpuid66] = 0;
            //check_bad_trap(spc66_phy_pc_w, 66, long_cpuid66);
            if(active_thread[long_cpuid66])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc66_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid66/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 66 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid66]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc66_phy_pc_w))
                begin
                    if(good[long_cpuid66/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid66 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid66/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid66])
        end // if (done[66])

        if (done[67]) begin
            timeout[long_cpuid67] = 0;
            //check_bad_trap(spc67_phy_pc_w, 67, long_cpuid67);
            if(active_thread[long_cpuid67])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc67_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid67/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 67 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid67]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc67_phy_pc_w))
                begin
                    if(good[long_cpuid67/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid67 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid67/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid67])
        end // if (done[67])

        if (done[68]) begin
            timeout[long_cpuid68] = 0;
            //check_bad_trap(spc68_phy_pc_w, 68, long_cpuid68);
            if(active_thread[long_cpuid68])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc68_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid68/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 68 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid68]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc68_phy_pc_w))
                begin
                    if(good[long_cpuid68/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid68 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid68/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid68])
        end // if (done[68])

        if (done[69]) begin
            timeout[long_cpuid69] = 0;
            //check_bad_trap(spc69_phy_pc_w, 69, long_cpuid69);
            if(active_thread[long_cpuid69])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc69_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid69/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 69 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid69]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc69_phy_pc_w))
                begin
                    if(good[long_cpuid69/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid69 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid69/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid69])
        end // if (done[69])

        if (done[70]) begin
            timeout[long_cpuid70] = 0;
            //check_bad_trap(spc70_phy_pc_w, 70, long_cpuid70);
            if(active_thread[long_cpuid70])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc70_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid70/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 70 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid70]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc70_phy_pc_w))
                begin
                    if(good[long_cpuid70/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid70 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid70/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid70])
        end // if (done[70])

        if (done[71]) begin
            timeout[long_cpuid71] = 0;
            //check_bad_trap(spc71_phy_pc_w, 71, long_cpuid71);
            if(active_thread[long_cpuid71])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc71_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid71/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 71 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid71]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc71_phy_pc_w))
                begin
                    if(good[long_cpuid71/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid71 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid71/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid71])
        end // if (done[71])

        if (done[72]) begin
            timeout[long_cpuid72] = 0;
            //check_bad_trap(spc72_phy_pc_w, 72, long_cpuid72);
            if(active_thread[long_cpuid72])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc72_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid72/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 72 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid72]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc72_phy_pc_w))
                begin
                    if(good[long_cpuid72/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid72 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid72/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid72])
        end // if (done[72])

        if (done[73]) begin
            timeout[long_cpuid73] = 0;
            //check_bad_trap(spc73_phy_pc_w, 73, long_cpuid73);
            if(active_thread[long_cpuid73])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc73_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid73/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 73 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid73]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc73_phy_pc_w))
                begin
                    if(good[long_cpuid73/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid73 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid73/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid73])
        end // if (done[73])

        if (done[74]) begin
            timeout[long_cpuid74] = 0;
            //check_bad_trap(spc74_phy_pc_w, 74, long_cpuid74);
            if(active_thread[long_cpuid74])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc74_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid74/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 74 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid74]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc74_phy_pc_w))
                begin
                    if(good[long_cpuid74/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid74 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid74/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid74])
        end // if (done[74])

        if (done[75]) begin
            timeout[long_cpuid75] = 0;
            //check_bad_trap(spc75_phy_pc_w, 75, long_cpuid75);
            if(active_thread[long_cpuid75])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc75_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid75/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 75 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid75]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc75_phy_pc_w))
                begin
                    if(good[long_cpuid75/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid75 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid75/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid75])
        end // if (done[75])

        if (done[76]) begin
            timeout[long_cpuid76] = 0;
            //check_bad_trap(spc76_phy_pc_w, 76, long_cpuid76);
            if(active_thread[long_cpuid76])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc76_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid76/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 76 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid76]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc76_phy_pc_w))
                begin
                    if(good[long_cpuid76/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid76 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid76/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid76])
        end // if (done[76])

        if (done[77]) begin
            timeout[long_cpuid77] = 0;
            //check_bad_trap(spc77_phy_pc_w, 77, long_cpuid77);
            if(active_thread[long_cpuid77])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc77_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid77/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 77 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid77]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc77_phy_pc_w))
                begin
                    if(good[long_cpuid77/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid77 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid77/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid77])
        end // if (done[77])

        if (done[78]) begin
            timeout[long_cpuid78] = 0;
            //check_bad_trap(spc78_phy_pc_w, 78, long_cpuid78);
            if(active_thread[long_cpuid78])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc78_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid78/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 78 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid78]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc78_phy_pc_w))
                begin
                    if(good[long_cpuid78/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid78 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid78/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid78])
        end // if (done[78])

        if (done[79]) begin
            timeout[long_cpuid79] = 0;
            //check_bad_trap(spc79_phy_pc_w, 79, long_cpuid79);
            if(active_thread[long_cpuid79])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc79_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid79/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 79 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid79]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc79_phy_pc_w))
                begin
                    if(good[long_cpuid79/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid79 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid79/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid79])
        end // if (done[79])

        if (done[80]) begin
            timeout[long_cpuid80] = 0;
            //check_bad_trap(spc80_phy_pc_w, 80, long_cpuid80);
            if(active_thread[long_cpuid80])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc80_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid80/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 80 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid80]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc80_phy_pc_w))
                begin
                    if(good[long_cpuid80/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid80 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid80/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid80])
        end // if (done[80])

        if (done[81]) begin
            timeout[long_cpuid81] = 0;
            //check_bad_trap(spc81_phy_pc_w, 81, long_cpuid81);
            if(active_thread[long_cpuid81])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc81_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid81/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 81 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid81]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc81_phy_pc_w))
                begin
                    if(good[long_cpuid81/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid81 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid81/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid81])
        end // if (done[81])

        if (done[82]) begin
            timeout[long_cpuid82] = 0;
            //check_bad_trap(spc82_phy_pc_w, 82, long_cpuid82);
            if(active_thread[long_cpuid82])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc82_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid82/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 82 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid82]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc82_phy_pc_w))
                begin
                    if(good[long_cpuid82/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid82 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid82/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid82])
        end // if (done[82])

        if (done[83]) begin
            timeout[long_cpuid83] = 0;
            //check_bad_trap(spc83_phy_pc_w, 83, long_cpuid83);
            if(active_thread[long_cpuid83])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc83_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid83/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 83 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid83]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc83_phy_pc_w))
                begin
                    if(good[long_cpuid83/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid83 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid83/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid83])
        end // if (done[83])

        if (done[84]) begin
            timeout[long_cpuid84] = 0;
            //check_bad_trap(spc84_phy_pc_w, 84, long_cpuid84);
            if(active_thread[long_cpuid84])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc84_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid84/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 84 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid84]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc84_phy_pc_w))
                begin
                    if(good[long_cpuid84/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid84 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid84/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid84])
        end // if (done[84])

        if (done[85]) begin
            timeout[long_cpuid85] = 0;
            //check_bad_trap(spc85_phy_pc_w, 85, long_cpuid85);
            if(active_thread[long_cpuid85])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc85_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid85/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 85 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid85]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc85_phy_pc_w))
                begin
                    if(good[long_cpuid85/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid85 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid85/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid85])
        end // if (done[85])

        if (done[86]) begin
            timeout[long_cpuid86] = 0;
            //check_bad_trap(spc86_phy_pc_w, 86, long_cpuid86);
            if(active_thread[long_cpuid86])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc86_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid86/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 86 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid86]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc86_phy_pc_w))
                begin
                    if(good[long_cpuid86/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid86 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid86/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid86])
        end // if (done[86])

        if (done[87]) begin
            timeout[long_cpuid87] = 0;
            //check_bad_trap(spc87_phy_pc_w, 87, long_cpuid87);
            if(active_thread[long_cpuid87])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc87_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid87/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 87 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid87]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc87_phy_pc_w))
                begin
                    if(good[long_cpuid87/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid87 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid87/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid87])
        end // if (done[87])

        if (done[88]) begin
            timeout[long_cpuid88] = 0;
            //check_bad_trap(spc88_phy_pc_w, 88, long_cpuid88);
            if(active_thread[long_cpuid88])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc88_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid88/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 88 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid88]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc88_phy_pc_w))
                begin
                    if(good[long_cpuid88/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid88 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid88/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid88])
        end // if (done[88])

        if (done[89]) begin
            timeout[long_cpuid89] = 0;
            //check_bad_trap(spc89_phy_pc_w, 89, long_cpuid89);
            if(active_thread[long_cpuid89])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc89_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid89/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 89 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid89]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc89_phy_pc_w))
                begin
                    if(good[long_cpuid89/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid89 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid89/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid89])
        end // if (done[89])

        if (done[90]) begin
            timeout[long_cpuid90] = 0;
            //check_bad_trap(spc90_phy_pc_w, 90, long_cpuid90);
            if(active_thread[long_cpuid90])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc90_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid90/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 90 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid90]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc90_phy_pc_w))
                begin
                    if(good[long_cpuid90/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid90 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid90/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid90])
        end // if (done[90])

        if (done[91]) begin
            timeout[long_cpuid91] = 0;
            //check_bad_trap(spc91_phy_pc_w, 91, long_cpuid91);
            if(active_thread[long_cpuid91])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc91_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid91/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 91 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid91]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc91_phy_pc_w))
                begin
                    if(good[long_cpuid91/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid91 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid91/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid91])
        end // if (done[91])

        if (done[92]) begin
            timeout[long_cpuid92] = 0;
            //check_bad_trap(spc92_phy_pc_w, 92, long_cpuid92);
            if(active_thread[long_cpuid92])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc92_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid92/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 92 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid92]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc92_phy_pc_w))
                begin
                    if(good[long_cpuid92/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid92 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid92/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid92])
        end // if (done[92])

        if (done[93]) begin
            timeout[long_cpuid93] = 0;
            //check_bad_trap(spc93_phy_pc_w, 93, long_cpuid93);
            if(active_thread[long_cpuid93])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc93_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid93/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 93 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid93]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc93_phy_pc_w))
                begin
                    if(good[long_cpuid93/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid93 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid93/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid93])
        end // if (done[93])

        if (done[94]) begin
            timeout[long_cpuid94] = 0;
            //check_bad_trap(spc94_phy_pc_w, 94, long_cpuid94);
            if(active_thread[long_cpuid94])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc94_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid94/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 94 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid94]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc94_phy_pc_w))
                begin
                    if(good[long_cpuid94/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid94 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid94/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid94])
        end // if (done[94])

        if (done[95]) begin
            timeout[long_cpuid95] = 0;
            //check_bad_trap(spc95_phy_pc_w, 95, long_cpuid95);
            if(active_thread[long_cpuid95])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc95_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid95/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 95 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid95]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc95_phy_pc_w))
                begin
                    if(good[long_cpuid95/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid95 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid95/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid95])
        end // if (done[95])

        if (done[96]) begin
            timeout[long_cpuid96] = 0;
            //check_bad_trap(spc96_phy_pc_w, 96, long_cpuid96);
            if(active_thread[long_cpuid96])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc96_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid96/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 96 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid96]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc96_phy_pc_w))
                begin
                    if(good[long_cpuid96/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid96 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid96/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid96])
        end // if (done[96])

        if (done[97]) begin
            timeout[long_cpuid97] = 0;
            //check_bad_trap(spc97_phy_pc_w, 97, long_cpuid97);
            if(active_thread[long_cpuid97])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc97_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid97/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 97 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid97]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc97_phy_pc_w))
                begin
                    if(good[long_cpuid97/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid97 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid97/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid97])
        end // if (done[97])

        if (done[98]) begin
            timeout[long_cpuid98] = 0;
            //check_bad_trap(spc98_phy_pc_w, 98, long_cpuid98);
            if(active_thread[long_cpuid98])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc98_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid98/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 98 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid98]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc98_phy_pc_w))
                begin
                    if(good[long_cpuid98/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid98 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid98/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid98])
        end // if (done[98])

        if (done[99]) begin
            timeout[long_cpuid99] = 0;
            //check_bad_trap(spc99_phy_pc_w, 99, long_cpuid99);
            if(active_thread[long_cpuid99])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc99_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid99/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 99 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid99]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc99_phy_pc_w))
                begin
                    if(good[long_cpuid99/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid99 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid99/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid99])
        end // if (done[99])

        if (done[100]) begin
            timeout[long_cpuid100] = 0;
            //check_bad_trap(spc100_phy_pc_w, 100, long_cpuid100);
            if(active_thread[long_cpuid100])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc100_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid100/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 100 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid100]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc100_phy_pc_w))
                begin
                    if(good[long_cpuid100/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid100 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid100/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid100])
        end // if (done[100])

        if (done[101]) begin
            timeout[long_cpuid101] = 0;
            //check_bad_trap(spc101_phy_pc_w, 101, long_cpuid101);
            if(active_thread[long_cpuid101])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc101_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid101/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 101 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid101]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc101_phy_pc_w))
                begin
                    if(good[long_cpuid101/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid101 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid101/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid101])
        end // if (done[101])

        if (done[102]) begin
            timeout[long_cpuid102] = 0;
            //check_bad_trap(spc102_phy_pc_w, 102, long_cpuid102);
            if(active_thread[long_cpuid102])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc102_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid102/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 102 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid102]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc102_phy_pc_w))
                begin
                    if(good[long_cpuid102/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid102 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid102/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid102])
        end // if (done[102])

        if (done[103]) begin
            timeout[long_cpuid103] = 0;
            //check_bad_trap(spc103_phy_pc_w, 103, long_cpuid103);
            if(active_thread[long_cpuid103])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc103_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid103/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 103 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid103]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc103_phy_pc_w))
                begin
                    if(good[long_cpuid103/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid103 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid103/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid103])
        end // if (done[103])

        if (done[104]) begin
            timeout[long_cpuid104] = 0;
            //check_bad_trap(spc104_phy_pc_w, 104, long_cpuid104);
            if(active_thread[long_cpuid104])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc104_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid104/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 104 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid104]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc104_phy_pc_w))
                begin
                    if(good[long_cpuid104/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid104 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid104/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid104])
        end // if (done[104])

        if (done[105]) begin
            timeout[long_cpuid105] = 0;
            //check_bad_trap(spc105_phy_pc_w, 105, long_cpuid105);
            if(active_thread[long_cpuid105])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc105_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid105/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 105 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid105]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc105_phy_pc_w))
                begin
                    if(good[long_cpuid105/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid105 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid105/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid105])
        end // if (done[105])

        if (done[106]) begin
            timeout[long_cpuid106] = 0;
            //check_bad_trap(spc106_phy_pc_w, 106, long_cpuid106);
            if(active_thread[long_cpuid106])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc106_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid106/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 106 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid106]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc106_phy_pc_w))
                begin
                    if(good[long_cpuid106/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid106 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid106/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid106])
        end // if (done[106])

        if (done[107]) begin
            timeout[long_cpuid107] = 0;
            //check_bad_trap(spc107_phy_pc_w, 107, long_cpuid107);
            if(active_thread[long_cpuid107])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc107_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid107/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 107 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid107]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc107_phy_pc_w))
                begin
                    if(good[long_cpuid107/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid107 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid107/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid107])
        end // if (done[107])

        if (done[108]) begin
            timeout[long_cpuid108] = 0;
            //check_bad_trap(spc108_phy_pc_w, 108, long_cpuid108);
            if(active_thread[long_cpuid108])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc108_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid108/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 108 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid108]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc108_phy_pc_w))
                begin
                    if(good[long_cpuid108/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid108 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid108/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid108])
        end // if (done[108])

        if (done[109]) begin
            timeout[long_cpuid109] = 0;
            //check_bad_trap(spc109_phy_pc_w, 109, long_cpuid109);
            if(active_thread[long_cpuid109])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc109_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid109/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 109 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid109]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc109_phy_pc_w))
                begin
                    if(good[long_cpuid109/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid109 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid109/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid109])
        end // if (done[109])

        if (done[110]) begin
            timeout[long_cpuid110] = 0;
            //check_bad_trap(spc110_phy_pc_w, 110, long_cpuid110);
            if(active_thread[long_cpuid110])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc110_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid110/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 110 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid110]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc110_phy_pc_w))
                begin
                    if(good[long_cpuid110/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid110 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid110/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid110])
        end // if (done[110])

        if (done[111]) begin
            timeout[long_cpuid111] = 0;
            //check_bad_trap(spc111_phy_pc_w, 111, long_cpuid111);
            if(active_thread[long_cpuid111])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc111_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid111/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 111 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid111]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc111_phy_pc_w))
                begin
                    if(good[long_cpuid111/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid111 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid111/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid111])
        end // if (done[111])

        if (done[112]) begin
            timeout[long_cpuid112] = 0;
            //check_bad_trap(spc112_phy_pc_w, 112, long_cpuid112);
            if(active_thread[long_cpuid112])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc112_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid112/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 112 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid112]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc112_phy_pc_w))
                begin
                    if(good[long_cpuid112/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid112 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid112/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid112])
        end // if (done[112])

        if (done[113]) begin
            timeout[long_cpuid113] = 0;
            //check_bad_trap(spc113_phy_pc_w, 113, long_cpuid113);
            if(active_thread[long_cpuid113])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc113_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid113/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 113 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid113]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc113_phy_pc_w))
                begin
                    if(good[long_cpuid113/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid113 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid113/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid113])
        end // if (done[113])

        if (done[114]) begin
            timeout[long_cpuid114] = 0;
            //check_bad_trap(spc114_phy_pc_w, 114, long_cpuid114);
            if(active_thread[long_cpuid114])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc114_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid114/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 114 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid114]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc114_phy_pc_w))
                begin
                    if(good[long_cpuid114/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid114 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid114/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid114])
        end // if (done[114])

        if (done[115]) begin
            timeout[long_cpuid115] = 0;
            //check_bad_trap(spc115_phy_pc_w, 115, long_cpuid115);
            if(active_thread[long_cpuid115])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc115_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid115/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 115 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid115]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc115_phy_pc_w))
                begin
                    if(good[long_cpuid115/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid115 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid115/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid115])
        end // if (done[115])

        if (done[116]) begin
            timeout[long_cpuid116] = 0;
            //check_bad_trap(spc116_phy_pc_w, 116, long_cpuid116);
            if(active_thread[long_cpuid116])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc116_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid116/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 116 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid116]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc116_phy_pc_w))
                begin
                    if(good[long_cpuid116/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid116 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid116/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid116])
        end // if (done[116])

        if (done[117]) begin
            timeout[long_cpuid117] = 0;
            //check_bad_trap(spc117_phy_pc_w, 117, long_cpuid117);
            if(active_thread[long_cpuid117])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc117_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid117/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 117 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid117]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc117_phy_pc_w))
                begin
                    if(good[long_cpuid117/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid117 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid117/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid117])
        end // if (done[117])

        if (done[118]) begin
            timeout[long_cpuid118] = 0;
            //check_bad_trap(spc118_phy_pc_w, 118, long_cpuid118);
            if(active_thread[long_cpuid118])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc118_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid118/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 118 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid118]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc118_phy_pc_w))
                begin
                    if(good[long_cpuid118/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid118 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid118/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid118])
        end // if (done[118])

        if (done[119]) begin
            timeout[long_cpuid119] = 0;
            //check_bad_trap(spc119_phy_pc_w, 119, long_cpuid119);
            if(active_thread[long_cpuid119])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc119_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid119/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 119 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid119]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc119_phy_pc_w))
                begin
                    if(good[long_cpuid119/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid119 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid119/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid119])
        end // if (done[119])

        if (done[120]) begin
            timeout[long_cpuid120] = 0;
            //check_bad_trap(spc120_phy_pc_w, 120, long_cpuid120);
            if(active_thread[long_cpuid120])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc120_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid120/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 120 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid120]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc120_phy_pc_w))
                begin
                    if(good[long_cpuid120/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid120 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid120/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid120])
        end // if (done[120])

        if (done[121]) begin
            timeout[long_cpuid121] = 0;
            //check_bad_trap(spc121_phy_pc_w, 121, long_cpuid121);
            if(active_thread[long_cpuid121])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc121_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid121/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 121 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid121]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc121_phy_pc_w))
                begin
                    if(good[long_cpuid121/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid121 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid121/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid121])
        end // if (done[121])

        if (done[122]) begin
            timeout[long_cpuid122] = 0;
            //check_bad_trap(spc122_phy_pc_w, 122, long_cpuid122);
            if(active_thread[long_cpuid122])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc122_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid122/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 122 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid122]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc122_phy_pc_w))
                begin
                    if(good[long_cpuid122/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid122 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid122/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid122])
        end // if (done[122])

        if (done[123]) begin
            timeout[long_cpuid123] = 0;
            //check_bad_trap(spc123_phy_pc_w, 123, long_cpuid123);
            if(active_thread[long_cpuid123])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc123_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid123/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 123 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid123]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc123_phy_pc_w))
                begin
                    if(good[long_cpuid123/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid123 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid123/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid123])
        end // if (done[123])

        if (done[124]) begin
            timeout[long_cpuid124] = 0;
            //check_bad_trap(spc124_phy_pc_w, 124, long_cpuid124);
            if(active_thread[long_cpuid124])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc124_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid124/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 124 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid124]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc124_phy_pc_w))
                begin
                    if(good[long_cpuid124/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid124 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid124/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid124])
        end // if (done[124])

        if (done[125]) begin
            timeout[long_cpuid125] = 0;
            //check_bad_trap(spc125_phy_pc_w, 125, long_cpuid125);
            if(active_thread[long_cpuid125])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc125_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid125/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 125 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid125]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc125_phy_pc_w))
                begin
                    if(good[long_cpuid125/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid125 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid125/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid125])
        end // if (done[125])

        if (done[126]) begin
            timeout[long_cpuid126] = 0;
            //check_bad_trap(spc126_phy_pc_w, 126, long_cpuid126);
            if(active_thread[long_cpuid126])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc126_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid126/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 126 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid126]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc126_phy_pc_w))
                begin
                    if(good[long_cpuid126/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid126 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid126/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid126])
        end // if (done[126])

        if (done[127]) begin
            timeout[long_cpuid127] = 0;
            //check_bad_trap(spc127_phy_pc_w, 127, long_cpuid127);
            if(active_thread[long_cpuid127])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc127_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid127/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 127 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid127]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc127_phy_pc_w))
                begin
                    if(good[long_cpuid127/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid127 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid127/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid127])
        end // if (done[127])

        if (done[128]) begin
            timeout[long_cpuid128] = 0;
            //check_bad_trap(spc128_phy_pc_w, 128, long_cpuid128);
            if(active_thread[long_cpuid128])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc128_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid128/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 128 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid128]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc128_phy_pc_w))
                begin
                    if(good[long_cpuid128/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid128 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid128/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid128])
        end // if (done[128])

        if (done[129]) begin
            timeout[long_cpuid129] = 0;
            //check_bad_trap(spc129_phy_pc_w, 129, long_cpuid129);
            if(active_thread[long_cpuid129])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc129_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid129/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 129 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid129]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc129_phy_pc_w))
                begin
                    if(good[long_cpuid129/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid129 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid129/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid129])
        end // if (done[129])

        if (done[130]) begin
            timeout[long_cpuid130] = 0;
            //check_bad_trap(spc130_phy_pc_w, 130, long_cpuid130);
            if(active_thread[long_cpuid130])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc130_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid130/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 130 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid130]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc130_phy_pc_w))
                begin
                    if(good[long_cpuid130/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid130 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid130/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid130])
        end // if (done[130])

        if (done[131]) begin
            timeout[long_cpuid131] = 0;
            //check_bad_trap(spc131_phy_pc_w, 131, long_cpuid131);
            if(active_thread[long_cpuid131])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc131_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid131/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 131 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid131]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc131_phy_pc_w))
                begin
                    if(good[long_cpuid131/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid131 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid131/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid131])
        end // if (done[131])

        if (done[132]) begin
            timeout[long_cpuid132] = 0;
            //check_bad_trap(spc132_phy_pc_w, 132, long_cpuid132);
            if(active_thread[long_cpuid132])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc132_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid132/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 132 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid132]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc132_phy_pc_w))
                begin
                    if(good[long_cpuid132/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid132 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid132/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid132])
        end // if (done[132])

        if (done[133]) begin
            timeout[long_cpuid133] = 0;
            //check_bad_trap(spc133_phy_pc_w, 133, long_cpuid133);
            if(active_thread[long_cpuid133])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc133_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid133/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 133 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid133]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc133_phy_pc_w))
                begin
                    if(good[long_cpuid133/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid133 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid133/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid133])
        end // if (done[133])

        if (done[134]) begin
            timeout[long_cpuid134] = 0;
            //check_bad_trap(spc134_phy_pc_w, 134, long_cpuid134);
            if(active_thread[long_cpuid134])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc134_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid134/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 134 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid134]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc134_phy_pc_w))
                begin
                    if(good[long_cpuid134/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid134 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid134/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid134])
        end // if (done[134])

        if (done[135]) begin
            timeout[long_cpuid135] = 0;
            //check_bad_trap(spc135_phy_pc_w, 135, long_cpuid135);
            if(active_thread[long_cpuid135])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc135_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid135/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 135 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid135]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc135_phy_pc_w))
                begin
                    if(good[long_cpuid135/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid135 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid135/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid135])
        end // if (done[135])

        if (done[136]) begin
            timeout[long_cpuid136] = 0;
            //check_bad_trap(spc136_phy_pc_w, 136, long_cpuid136);
            if(active_thread[long_cpuid136])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc136_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid136/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 136 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid136]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc136_phy_pc_w))
                begin
                    if(good[long_cpuid136/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid136 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid136/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid136])
        end // if (done[136])

        if (done[137]) begin
            timeout[long_cpuid137] = 0;
            //check_bad_trap(spc137_phy_pc_w, 137, long_cpuid137);
            if(active_thread[long_cpuid137])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc137_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid137/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 137 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid137]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc137_phy_pc_w))
                begin
                    if(good[long_cpuid137/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid137 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid137/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid137])
        end // if (done[137])

        if (done[138]) begin
            timeout[long_cpuid138] = 0;
            //check_bad_trap(spc138_phy_pc_w, 138, long_cpuid138);
            if(active_thread[long_cpuid138])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc138_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid138/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 138 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid138]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc138_phy_pc_w))
                begin
                    if(good[long_cpuid138/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid138 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid138/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid138])
        end // if (done[138])

        if (done[139]) begin
            timeout[long_cpuid139] = 0;
            //check_bad_trap(spc139_phy_pc_w, 139, long_cpuid139);
            if(active_thread[long_cpuid139])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc139_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid139/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 139 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid139]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc139_phy_pc_w))
                begin
                    if(good[long_cpuid139/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid139 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid139/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid139])
        end // if (done[139])

        if (done[140]) begin
            timeout[long_cpuid140] = 0;
            //check_bad_trap(spc140_phy_pc_w, 140, long_cpuid140);
            if(active_thread[long_cpuid140])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc140_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid140/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 140 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid140]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc140_phy_pc_w))
                begin
                    if(good[long_cpuid140/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid140 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid140/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid140])
        end // if (done[140])

        if (done[141]) begin
            timeout[long_cpuid141] = 0;
            //check_bad_trap(spc141_phy_pc_w, 141, long_cpuid141);
            if(active_thread[long_cpuid141])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc141_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid141/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 141 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid141]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc141_phy_pc_w))
                begin
                    if(good[long_cpuid141/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid141 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid141/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid141])
        end // if (done[141])

        if (done[142]) begin
            timeout[long_cpuid142] = 0;
            //check_bad_trap(spc142_phy_pc_w, 142, long_cpuid142);
            if(active_thread[long_cpuid142])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc142_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid142/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 142 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid142]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc142_phy_pc_w))
                begin
                    if(good[long_cpuid142/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid142 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid142/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid142])
        end // if (done[142])

        if (done[143]) begin
            timeout[long_cpuid143] = 0;
            //check_bad_trap(spc143_phy_pc_w, 143, long_cpuid143);
            if(active_thread[long_cpuid143])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc143_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid143/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 143 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid143]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc143_phy_pc_w))
                begin
                    if(good[long_cpuid143/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid143 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid143/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid143])
        end // if (done[143])

        if (done[144]) begin
            timeout[long_cpuid144] = 0;
            //check_bad_trap(spc144_phy_pc_w, 144, long_cpuid144);
            if(active_thread[long_cpuid144])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc144_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid144/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 144 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid144]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc144_phy_pc_w))
                begin
                    if(good[long_cpuid144/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid144 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid144/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid144])
        end // if (done[144])

        if (done[145]) begin
            timeout[long_cpuid145] = 0;
            //check_bad_trap(spc145_phy_pc_w, 145, long_cpuid145);
            if(active_thread[long_cpuid145])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc145_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid145/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 145 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid145]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc145_phy_pc_w))
                begin
                    if(good[long_cpuid145/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid145 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid145/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid145])
        end // if (done[145])

        if (done[146]) begin
            timeout[long_cpuid146] = 0;
            //check_bad_trap(spc146_phy_pc_w, 146, long_cpuid146);
            if(active_thread[long_cpuid146])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc146_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid146/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 146 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid146]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc146_phy_pc_w))
                begin
                    if(good[long_cpuid146/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid146 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid146/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid146])
        end // if (done[146])

        if (done[147]) begin
            timeout[long_cpuid147] = 0;
            //check_bad_trap(spc147_phy_pc_w, 147, long_cpuid147);
            if(active_thread[long_cpuid147])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc147_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid147/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 147 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid147]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc147_phy_pc_w))
                begin
                    if(good[long_cpuid147/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid147 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid147/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid147])
        end // if (done[147])

        if (done[148]) begin
            timeout[long_cpuid148] = 0;
            //check_bad_trap(spc148_phy_pc_w, 148, long_cpuid148);
            if(active_thread[long_cpuid148])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc148_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid148/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 148 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid148]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc148_phy_pc_w))
                begin
                    if(good[long_cpuid148/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid148 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid148/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid148])
        end // if (done[148])

        if (done[149]) begin
            timeout[long_cpuid149] = 0;
            //check_bad_trap(spc149_phy_pc_w, 149, long_cpuid149);
            if(active_thread[long_cpuid149])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc149_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid149/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 149 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid149]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc149_phy_pc_w))
                begin
                    if(good[long_cpuid149/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid149 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid149/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid149])
        end // if (done[149])

        if (done[150]) begin
            timeout[long_cpuid150] = 0;
            //check_bad_trap(spc150_phy_pc_w, 150, long_cpuid150);
            if(active_thread[long_cpuid150])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc150_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid150/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 150 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid150]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc150_phy_pc_w))
                begin
                    if(good[long_cpuid150/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid150 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid150/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid150])
        end // if (done[150])

        if (done[151]) begin
            timeout[long_cpuid151] = 0;
            //check_bad_trap(spc151_phy_pc_w, 151, long_cpuid151);
            if(active_thread[long_cpuid151])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc151_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid151/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 151 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid151]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc151_phy_pc_w))
                begin
                    if(good[long_cpuid151/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid151 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid151/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid151])
        end // if (done[151])

        if (done[152]) begin
            timeout[long_cpuid152] = 0;
            //check_bad_trap(spc152_phy_pc_w, 152, long_cpuid152);
            if(active_thread[long_cpuid152])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc152_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid152/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 152 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid152]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc152_phy_pc_w))
                begin
                    if(good[long_cpuid152/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid152 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid152/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid152])
        end // if (done[152])

        if (done[153]) begin
            timeout[long_cpuid153] = 0;
            //check_bad_trap(spc153_phy_pc_w, 153, long_cpuid153);
            if(active_thread[long_cpuid153])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc153_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid153/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 153 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid153]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc153_phy_pc_w))
                begin
                    if(good[long_cpuid153/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid153 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid153/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid153])
        end // if (done[153])

        if (done[154]) begin
            timeout[long_cpuid154] = 0;
            //check_bad_trap(spc154_phy_pc_w, 154, long_cpuid154);
            if(active_thread[long_cpuid154])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc154_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid154/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 154 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid154]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc154_phy_pc_w))
                begin
                    if(good[long_cpuid154/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid154 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid154/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid154])
        end // if (done[154])

        if (done[155]) begin
            timeout[long_cpuid155] = 0;
            //check_bad_trap(spc155_phy_pc_w, 155, long_cpuid155);
            if(active_thread[long_cpuid155])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc155_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid155/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 155 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid155]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc155_phy_pc_w))
                begin
                    if(good[long_cpuid155/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid155 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid155/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid155])
        end // if (done[155])

        if (done[156]) begin
            timeout[long_cpuid156] = 0;
            //check_bad_trap(spc156_phy_pc_w, 156, long_cpuid156);
            if(active_thread[long_cpuid156])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc156_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid156/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 156 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid156]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc156_phy_pc_w))
                begin
                    if(good[long_cpuid156/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid156 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid156/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid156])
        end // if (done[156])

        if (done[157]) begin
            timeout[long_cpuid157] = 0;
            //check_bad_trap(spc157_phy_pc_w, 157, long_cpuid157);
            if(active_thread[long_cpuid157])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc157_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid157/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 157 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid157]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc157_phy_pc_w))
                begin
                    if(good[long_cpuid157/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid157 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid157/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid157])
        end // if (done[157])

        if (done[158]) begin
            timeout[long_cpuid158] = 0;
            //check_bad_trap(spc158_phy_pc_w, 158, long_cpuid158);
            if(active_thread[long_cpuid158])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc158_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid158/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 158 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid158]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc158_phy_pc_w))
                begin
                    if(good[long_cpuid158/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid158 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid158/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid158])
        end // if (done[158])

        if (done[159]) begin
            timeout[long_cpuid159] = 0;
            //check_bad_trap(spc159_phy_pc_w, 159, long_cpuid159);
            if(active_thread[long_cpuid159])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc159_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid159/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 159 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid159]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc159_phy_pc_w))
                begin
                    if(good[long_cpuid159/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid159 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid159/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid159])
        end // if (done[159])

        if (done[160]) begin
            timeout[long_cpuid160] = 0;
            //check_bad_trap(spc160_phy_pc_w, 160, long_cpuid160);
            if(active_thread[long_cpuid160])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc160_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid160/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 160 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid160]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc160_phy_pc_w))
                begin
                    if(good[long_cpuid160/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid160 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid160/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid160])
        end // if (done[160])

        if (done[161]) begin
            timeout[long_cpuid161] = 0;
            //check_bad_trap(spc161_phy_pc_w, 161, long_cpuid161);
            if(active_thread[long_cpuid161])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc161_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid161/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 161 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid161]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc161_phy_pc_w))
                begin
                    if(good[long_cpuid161/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid161 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid161/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid161])
        end // if (done[161])

        if (done[162]) begin
            timeout[long_cpuid162] = 0;
            //check_bad_trap(spc162_phy_pc_w, 162, long_cpuid162);
            if(active_thread[long_cpuid162])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc162_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid162/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 162 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid162]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc162_phy_pc_w))
                begin
                    if(good[long_cpuid162/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid162 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid162/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid162])
        end // if (done[162])

        if (done[163]) begin
            timeout[long_cpuid163] = 0;
            //check_bad_trap(spc163_phy_pc_w, 163, long_cpuid163);
            if(active_thread[long_cpuid163])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc163_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid163/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 163 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid163]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc163_phy_pc_w))
                begin
                    if(good[long_cpuid163/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid163 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid163/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid163])
        end // if (done[163])

        if (done[164]) begin
            timeout[long_cpuid164] = 0;
            //check_bad_trap(spc164_phy_pc_w, 164, long_cpuid164);
            if(active_thread[long_cpuid164])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc164_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid164/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 164 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid164]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc164_phy_pc_w))
                begin
                    if(good[long_cpuid164/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid164 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid164/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid164])
        end // if (done[164])

        if (done[165]) begin
            timeout[long_cpuid165] = 0;
            //check_bad_trap(spc165_phy_pc_w, 165, long_cpuid165);
            if(active_thread[long_cpuid165])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc165_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid165/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 165 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid165]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc165_phy_pc_w))
                begin
                    if(good[long_cpuid165/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid165 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid165/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid165])
        end // if (done[165])

        if (done[166]) begin
            timeout[long_cpuid166] = 0;
            //check_bad_trap(spc166_phy_pc_w, 166, long_cpuid166);
            if(active_thread[long_cpuid166])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc166_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid166/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 166 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid166]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc166_phy_pc_w))
                begin
                    if(good[long_cpuid166/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid166 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid166/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid166])
        end // if (done[166])

        if (done[167]) begin
            timeout[long_cpuid167] = 0;
            //check_bad_trap(spc167_phy_pc_w, 167, long_cpuid167);
            if(active_thread[long_cpuid167])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc167_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid167/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 167 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid167]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc167_phy_pc_w))
                begin
                    if(good[long_cpuid167/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid167 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid167/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid167])
        end // if (done[167])

        if (done[168]) begin
            timeout[long_cpuid168] = 0;
            //check_bad_trap(spc168_phy_pc_w, 168, long_cpuid168);
            if(active_thread[long_cpuid168])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc168_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid168/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 168 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid168]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc168_phy_pc_w))
                begin
                    if(good[long_cpuid168/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid168 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid168/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid168])
        end // if (done[168])

        if (done[169]) begin
            timeout[long_cpuid169] = 0;
            //check_bad_trap(spc169_phy_pc_w, 169, long_cpuid169);
            if(active_thread[long_cpuid169])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc169_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid169/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 169 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid169]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc169_phy_pc_w))
                begin
                    if(good[long_cpuid169/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid169 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid169/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid169])
        end // if (done[169])

        if (done[170]) begin
            timeout[long_cpuid170] = 0;
            //check_bad_trap(spc170_phy_pc_w, 170, long_cpuid170);
            if(active_thread[long_cpuid170])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc170_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid170/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 170 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid170]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc170_phy_pc_w))
                begin
                    if(good[long_cpuid170/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid170 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid170/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid170])
        end // if (done[170])

        if (done[171]) begin
            timeout[long_cpuid171] = 0;
            //check_bad_trap(spc171_phy_pc_w, 171, long_cpuid171);
            if(active_thread[long_cpuid171])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc171_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid171/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 171 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid171]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc171_phy_pc_w))
                begin
                    if(good[long_cpuid171/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid171 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid171/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid171])
        end // if (done[171])

        if (done[172]) begin
            timeout[long_cpuid172] = 0;
            //check_bad_trap(spc172_phy_pc_w, 172, long_cpuid172);
            if(active_thread[long_cpuid172])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc172_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid172/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 172 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid172]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc172_phy_pc_w))
                begin
                    if(good[long_cpuid172/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid172 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid172/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid172])
        end // if (done[172])

        if (done[173]) begin
            timeout[long_cpuid173] = 0;
            //check_bad_trap(spc173_phy_pc_w, 173, long_cpuid173);
            if(active_thread[long_cpuid173])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc173_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid173/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 173 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid173]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc173_phy_pc_w))
                begin
                    if(good[long_cpuid173/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid173 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid173/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid173])
        end // if (done[173])

        if (done[174]) begin
            timeout[long_cpuid174] = 0;
            //check_bad_trap(spc174_phy_pc_w, 174, long_cpuid174);
            if(active_thread[long_cpuid174])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc174_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid174/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 174 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid174]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc174_phy_pc_w))
                begin
                    if(good[long_cpuid174/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid174 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid174/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid174])
        end // if (done[174])

        if (done[175]) begin
            timeout[long_cpuid175] = 0;
            //check_bad_trap(spc175_phy_pc_w, 175, long_cpuid175);
            if(active_thread[long_cpuid175])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc175_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid175/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 175 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid175]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc175_phy_pc_w))
                begin
                    if(good[long_cpuid175/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid175 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid175/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid175])
        end // if (done[175])

        if (done[176]) begin
            timeout[long_cpuid176] = 0;
            //check_bad_trap(spc176_phy_pc_w, 176, long_cpuid176);
            if(active_thread[long_cpuid176])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc176_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid176/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 176 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid176]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc176_phy_pc_w))
                begin
                    if(good[long_cpuid176/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid176 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid176/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid176])
        end // if (done[176])

        if (done[177]) begin
            timeout[long_cpuid177] = 0;
            //check_bad_trap(spc177_phy_pc_w, 177, long_cpuid177);
            if(active_thread[long_cpuid177])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc177_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid177/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 177 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid177]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc177_phy_pc_w))
                begin
                    if(good[long_cpuid177/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid177 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid177/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid177])
        end // if (done[177])

        if (done[178]) begin
            timeout[long_cpuid178] = 0;
            //check_bad_trap(spc178_phy_pc_w, 178, long_cpuid178);
            if(active_thread[long_cpuid178])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc178_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid178/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 178 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid178]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc178_phy_pc_w))
                begin
                    if(good[long_cpuid178/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid178 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid178/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid178])
        end // if (done[178])

        if (done[179]) begin
            timeout[long_cpuid179] = 0;
            //check_bad_trap(spc179_phy_pc_w, 179, long_cpuid179);
            if(active_thread[long_cpuid179])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc179_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid179/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 179 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid179]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc179_phy_pc_w))
                begin
                    if(good[long_cpuid179/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid179 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid179/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid179])
        end // if (done[179])

        if (done[180]) begin
            timeout[long_cpuid180] = 0;
            //check_bad_trap(spc180_phy_pc_w, 180, long_cpuid180);
            if(active_thread[long_cpuid180])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc180_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid180/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 180 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid180]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc180_phy_pc_w))
                begin
                    if(good[long_cpuid180/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid180 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid180/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid180])
        end // if (done[180])

        if (done[181]) begin
            timeout[long_cpuid181] = 0;
            //check_bad_trap(spc181_phy_pc_w, 181, long_cpuid181);
            if(active_thread[long_cpuid181])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc181_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid181/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 181 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid181]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc181_phy_pc_w))
                begin
                    if(good[long_cpuid181/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid181 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid181/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid181])
        end // if (done[181])

        if (done[182]) begin
            timeout[long_cpuid182] = 0;
            //check_bad_trap(spc182_phy_pc_w, 182, long_cpuid182);
            if(active_thread[long_cpuid182])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc182_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid182/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 182 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid182]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc182_phy_pc_w))
                begin
                    if(good[long_cpuid182/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid182 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid182/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid182])
        end // if (done[182])

        if (done[183]) begin
            timeout[long_cpuid183] = 0;
            //check_bad_trap(spc183_phy_pc_w, 183, long_cpuid183);
            if(active_thread[long_cpuid183])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc183_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid183/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 183 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid183]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc183_phy_pc_w))
                begin
                    if(good[long_cpuid183/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid183 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid183/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid183])
        end // if (done[183])

        if (done[184]) begin
            timeout[long_cpuid184] = 0;
            //check_bad_trap(spc184_phy_pc_w, 184, long_cpuid184);
            if(active_thread[long_cpuid184])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc184_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid184/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 184 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid184]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc184_phy_pc_w))
                begin
                    if(good[long_cpuid184/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid184 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid184/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid184])
        end // if (done[184])

        if (done[185]) begin
            timeout[long_cpuid185] = 0;
            //check_bad_trap(spc185_phy_pc_w, 185, long_cpuid185);
            if(active_thread[long_cpuid185])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc185_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid185/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 185 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid185]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc185_phy_pc_w))
                begin
                    if(good[long_cpuid185/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid185 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid185/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid185])
        end // if (done[185])

        if (done[186]) begin
            timeout[long_cpuid186] = 0;
            //check_bad_trap(spc186_phy_pc_w, 186, long_cpuid186);
            if(active_thread[long_cpuid186])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc186_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid186/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 186 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid186]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc186_phy_pc_w))
                begin
                    if(good[long_cpuid186/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid186 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid186/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid186])
        end // if (done[186])

        if (done[187]) begin
            timeout[long_cpuid187] = 0;
            //check_bad_trap(spc187_phy_pc_w, 187, long_cpuid187);
            if(active_thread[long_cpuid187])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc187_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid187/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 187 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid187]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc187_phy_pc_w))
                begin
                    if(good[long_cpuid187/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid187 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid187/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid187])
        end // if (done[187])

        if (done[188]) begin
            timeout[long_cpuid188] = 0;
            //check_bad_trap(spc188_phy_pc_w, 188, long_cpuid188);
            if(active_thread[long_cpuid188])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc188_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid188/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 188 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid188]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc188_phy_pc_w))
                begin
                    if(good[long_cpuid188/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid188 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid188/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid188])
        end // if (done[188])

        if (done[189]) begin
            timeout[long_cpuid189] = 0;
            //check_bad_trap(spc189_phy_pc_w, 189, long_cpuid189);
            if(active_thread[long_cpuid189])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc189_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid189/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 189 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid189]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc189_phy_pc_w))
                begin
                    if(good[long_cpuid189/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid189 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid189/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid189])
        end // if (done[189])

        if (done[190]) begin
            timeout[long_cpuid190] = 0;
            //check_bad_trap(spc190_phy_pc_w, 190, long_cpuid190);
            if(active_thread[long_cpuid190])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc190_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid190/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 190 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid190]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc190_phy_pc_w))
                begin
                    if(good[long_cpuid190/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid190 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid190/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid190])
        end // if (done[190])

        if (done[191]) begin
            timeout[long_cpuid191] = 0;
            //check_bad_trap(spc191_phy_pc_w, 191, long_cpuid191);
            if(active_thread[long_cpuid191])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc191_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid191/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 191 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid191]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc191_phy_pc_w))
                begin
                    if(good[long_cpuid191/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid191 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid191/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid191])
        end // if (done[191])

        if (done[192]) begin
            timeout[long_cpuid192] = 0;
            //check_bad_trap(spc192_phy_pc_w, 192, long_cpuid192);
            if(active_thread[long_cpuid192])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc192_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid192/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 192 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid192]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc192_phy_pc_w))
                begin
                    if(good[long_cpuid192/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid192 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid192/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid192])
        end // if (done[192])

        if (done[193]) begin
            timeout[long_cpuid193] = 0;
            //check_bad_trap(spc193_phy_pc_w, 193, long_cpuid193);
            if(active_thread[long_cpuid193])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc193_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid193/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 193 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid193]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc193_phy_pc_w))
                begin
                    if(good[long_cpuid193/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid193 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid193/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid193])
        end // if (done[193])

        if (done[194]) begin
            timeout[long_cpuid194] = 0;
            //check_bad_trap(spc194_phy_pc_w, 194, long_cpuid194);
            if(active_thread[long_cpuid194])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc194_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid194/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 194 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid194]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc194_phy_pc_w))
                begin
                    if(good[long_cpuid194/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid194 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid194/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid194])
        end // if (done[194])

        if (done[195]) begin
            timeout[long_cpuid195] = 0;
            //check_bad_trap(spc195_phy_pc_w, 195, long_cpuid195);
            if(active_thread[long_cpuid195])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc195_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid195/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 195 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid195]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc195_phy_pc_w))
                begin
                    if(good[long_cpuid195/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid195 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid195/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid195])
        end // if (done[195])

        if (done[196]) begin
            timeout[long_cpuid196] = 0;
            //check_bad_trap(spc196_phy_pc_w, 196, long_cpuid196);
            if(active_thread[long_cpuid196])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc196_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid196/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 196 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid196]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc196_phy_pc_w))
                begin
                    if(good[long_cpuid196/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid196 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid196/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid196])
        end // if (done[196])

        if (done[197]) begin
            timeout[long_cpuid197] = 0;
            //check_bad_trap(spc197_phy_pc_w, 197, long_cpuid197);
            if(active_thread[long_cpuid197])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc197_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid197/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 197 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid197]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc197_phy_pc_w))
                begin
                    if(good[long_cpuid197/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid197 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid197/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid197])
        end // if (done[197])

        if (done[198]) begin
            timeout[long_cpuid198] = 0;
            //check_bad_trap(spc198_phy_pc_w, 198, long_cpuid198);
            if(active_thread[long_cpuid198])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc198_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid198/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 198 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid198]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc198_phy_pc_w))
                begin
                    if(good[long_cpuid198/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid198 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid198/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid198])
        end // if (done[198])

        if (done[199]) begin
            timeout[long_cpuid199] = 0;
            //check_bad_trap(spc199_phy_pc_w, 199, long_cpuid199);
            if(active_thread[long_cpuid199])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc199_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid199/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 199 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid199]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc199_phy_pc_w))
                begin
                    if(good[long_cpuid199/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid199 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid199/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid199])
        end // if (done[199])

        if (done[200]) begin
            timeout[long_cpuid200] = 0;
            //check_bad_trap(spc200_phy_pc_w, 200, long_cpuid200);
            if(active_thread[long_cpuid200])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc200_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid200/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 200 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid200]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc200_phy_pc_w))
                begin
                    if(good[long_cpuid200/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid200 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid200/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid200])
        end // if (done[200])

        if (done[201]) begin
            timeout[long_cpuid201] = 0;
            //check_bad_trap(spc201_phy_pc_w, 201, long_cpuid201);
            if(active_thread[long_cpuid201])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc201_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid201/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 201 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid201]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc201_phy_pc_w))
                begin
                    if(good[long_cpuid201/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid201 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid201/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid201])
        end // if (done[201])

        if (done[202]) begin
            timeout[long_cpuid202] = 0;
            //check_bad_trap(spc202_phy_pc_w, 202, long_cpuid202);
            if(active_thread[long_cpuid202])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc202_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid202/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 202 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid202]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc202_phy_pc_w))
                begin
                    if(good[long_cpuid202/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid202 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid202/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid202])
        end // if (done[202])

        if (done[203]) begin
            timeout[long_cpuid203] = 0;
            //check_bad_trap(spc203_phy_pc_w, 203, long_cpuid203);
            if(active_thread[long_cpuid203])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc203_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid203/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 203 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid203]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc203_phy_pc_w))
                begin
                    if(good[long_cpuid203/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid203 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid203/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid203])
        end // if (done[203])

        if (done[204]) begin
            timeout[long_cpuid204] = 0;
            //check_bad_trap(spc204_phy_pc_w, 204, long_cpuid204);
            if(active_thread[long_cpuid204])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc204_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid204/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 204 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid204]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc204_phy_pc_w))
                begin
                    if(good[long_cpuid204/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid204 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid204/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid204])
        end // if (done[204])

        if (done[205]) begin
            timeout[long_cpuid205] = 0;
            //check_bad_trap(spc205_phy_pc_w, 205, long_cpuid205);
            if(active_thread[long_cpuid205])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc205_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid205/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 205 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid205]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc205_phy_pc_w))
                begin
                    if(good[long_cpuid205/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid205 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid205/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid205])
        end // if (done[205])

        if (done[206]) begin
            timeout[long_cpuid206] = 0;
            //check_bad_trap(spc206_phy_pc_w, 206, long_cpuid206);
            if(active_thread[long_cpuid206])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc206_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid206/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 206 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid206]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc206_phy_pc_w))
                begin
                    if(good[long_cpuid206/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid206 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid206/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid206])
        end // if (done[206])

        if (done[207]) begin
            timeout[long_cpuid207] = 0;
            //check_bad_trap(spc207_phy_pc_w, 207, long_cpuid207);
            if(active_thread[long_cpuid207])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc207_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid207/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 207 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid207]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc207_phy_pc_w))
                begin
                    if(good[long_cpuid207/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid207 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid207/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid207])
        end // if (done[207])

        if (done[208]) begin
            timeout[long_cpuid208] = 0;
            //check_bad_trap(spc208_phy_pc_w, 208, long_cpuid208);
            if(active_thread[long_cpuid208])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc208_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid208/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 208 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid208]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc208_phy_pc_w))
                begin
                    if(good[long_cpuid208/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid208 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid208/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid208])
        end // if (done[208])

        if (done[209]) begin
            timeout[long_cpuid209] = 0;
            //check_bad_trap(spc209_phy_pc_w, 209, long_cpuid209);
            if(active_thread[long_cpuid209])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc209_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid209/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 209 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid209]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc209_phy_pc_w))
                begin
                    if(good[long_cpuid209/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid209 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid209/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid209])
        end // if (done[209])

        if (done[210]) begin
            timeout[long_cpuid210] = 0;
            //check_bad_trap(spc210_phy_pc_w, 210, long_cpuid210);
            if(active_thread[long_cpuid210])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc210_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid210/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 210 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid210]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc210_phy_pc_w))
                begin
                    if(good[long_cpuid210/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid210 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid210/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid210])
        end // if (done[210])

        if (done[211]) begin
            timeout[long_cpuid211] = 0;
            //check_bad_trap(spc211_phy_pc_w, 211, long_cpuid211);
            if(active_thread[long_cpuid211])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc211_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid211/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 211 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid211]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc211_phy_pc_w))
                begin
                    if(good[long_cpuid211/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid211 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid211/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid211])
        end // if (done[211])

        if (done[212]) begin
            timeout[long_cpuid212] = 0;
            //check_bad_trap(spc212_phy_pc_w, 212, long_cpuid212);
            if(active_thread[long_cpuid212])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc212_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid212/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 212 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid212]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc212_phy_pc_w))
                begin
                    if(good[long_cpuid212/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid212 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid212/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid212])
        end // if (done[212])

        if (done[213]) begin
            timeout[long_cpuid213] = 0;
            //check_bad_trap(spc213_phy_pc_w, 213, long_cpuid213);
            if(active_thread[long_cpuid213])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc213_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid213/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 213 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid213]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc213_phy_pc_w))
                begin
                    if(good[long_cpuid213/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid213 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid213/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid213])
        end // if (done[213])

        if (done[214]) begin
            timeout[long_cpuid214] = 0;
            //check_bad_trap(spc214_phy_pc_w, 214, long_cpuid214);
            if(active_thread[long_cpuid214])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc214_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid214/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 214 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid214]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc214_phy_pc_w))
                begin
                    if(good[long_cpuid214/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid214 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid214/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid214])
        end // if (done[214])

        if (done[215]) begin
            timeout[long_cpuid215] = 0;
            //check_bad_trap(spc215_phy_pc_w, 215, long_cpuid215);
            if(active_thread[long_cpuid215])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc215_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid215/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 215 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid215]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc215_phy_pc_w))
                begin
                    if(good[long_cpuid215/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid215 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid215/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid215])
        end // if (done[215])

        if (done[216]) begin
            timeout[long_cpuid216] = 0;
            //check_bad_trap(spc216_phy_pc_w, 216, long_cpuid216);
            if(active_thread[long_cpuid216])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc216_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid216/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 216 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid216]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc216_phy_pc_w))
                begin
                    if(good[long_cpuid216/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid216 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid216/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid216])
        end // if (done[216])

        if (done[217]) begin
            timeout[long_cpuid217] = 0;
            //check_bad_trap(spc217_phy_pc_w, 217, long_cpuid217);
            if(active_thread[long_cpuid217])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc217_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid217/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 217 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid217]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc217_phy_pc_w))
                begin
                    if(good[long_cpuid217/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid217 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid217/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid217])
        end // if (done[217])

        if (done[218]) begin
            timeout[long_cpuid218] = 0;
            //check_bad_trap(spc218_phy_pc_w, 218, long_cpuid218);
            if(active_thread[long_cpuid218])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc218_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid218/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 218 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid218]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc218_phy_pc_w))
                begin
                    if(good[long_cpuid218/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid218 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid218/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid218])
        end // if (done[218])

        if (done[219]) begin
            timeout[long_cpuid219] = 0;
            //check_bad_trap(spc219_phy_pc_w, 219, long_cpuid219);
            if(active_thread[long_cpuid219])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc219_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid219/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 219 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid219]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc219_phy_pc_w))
                begin
                    if(good[long_cpuid219/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid219 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid219/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid219])
        end // if (done[219])

        if (done[220]) begin
            timeout[long_cpuid220] = 0;
            //check_bad_trap(spc220_phy_pc_w, 220, long_cpuid220);
            if(active_thread[long_cpuid220])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc220_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid220/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 220 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid220]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc220_phy_pc_w))
                begin
                    if(good[long_cpuid220/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid220 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid220/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid220])
        end // if (done[220])

        if (done[221]) begin
            timeout[long_cpuid221] = 0;
            //check_bad_trap(spc221_phy_pc_w, 221, long_cpuid221);
            if(active_thread[long_cpuid221])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc221_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid221/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 221 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid221]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc221_phy_pc_w))
                begin
                    if(good[long_cpuid221/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid221 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid221/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid221])
        end // if (done[221])

        if (done[222]) begin
            timeout[long_cpuid222] = 0;
            //check_bad_trap(spc222_phy_pc_w, 222, long_cpuid222);
            if(active_thread[long_cpuid222])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc222_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid222/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 222 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid222]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc222_phy_pc_w))
                begin
                    if(good[long_cpuid222/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid222 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid222/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid222])
        end // if (done[222])

        if (done[223]) begin
            timeout[long_cpuid223] = 0;
            //check_bad_trap(spc223_phy_pc_w, 223, long_cpuid223);
            if(active_thread[long_cpuid223])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc223_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid223/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 223 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid223]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc223_phy_pc_w))
                begin
                    if(good[long_cpuid223/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid223 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid223/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid223])
        end // if (done[223])

        if (done[224]) begin
            timeout[long_cpuid224] = 0;
            //check_bad_trap(spc224_phy_pc_w, 224, long_cpuid224);
            if(active_thread[long_cpuid224])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc224_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid224/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 224 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid224]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc224_phy_pc_w))
                begin
                    if(good[long_cpuid224/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid224 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid224/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid224])
        end // if (done[224])

        if (done[225]) begin
            timeout[long_cpuid225] = 0;
            //check_bad_trap(spc225_phy_pc_w, 225, long_cpuid225);
            if(active_thread[long_cpuid225])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc225_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid225/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 225 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid225]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc225_phy_pc_w))
                begin
                    if(good[long_cpuid225/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid225 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid225/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid225])
        end // if (done[225])

        if (done[226]) begin
            timeout[long_cpuid226] = 0;
            //check_bad_trap(spc226_phy_pc_w, 226, long_cpuid226);
            if(active_thread[long_cpuid226])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc226_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid226/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 226 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid226]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc226_phy_pc_w))
                begin
                    if(good[long_cpuid226/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid226 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid226/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid226])
        end // if (done[226])

        if (done[227]) begin
            timeout[long_cpuid227] = 0;
            //check_bad_trap(spc227_phy_pc_w, 227, long_cpuid227);
            if(active_thread[long_cpuid227])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc227_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid227/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 227 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid227]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc227_phy_pc_w))
                begin
                    if(good[long_cpuid227/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid227 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid227/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid227])
        end // if (done[227])

        if (done[228]) begin
            timeout[long_cpuid228] = 0;
            //check_bad_trap(spc228_phy_pc_w, 228, long_cpuid228);
            if(active_thread[long_cpuid228])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc228_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid228/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 228 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid228]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc228_phy_pc_w))
                begin
                    if(good[long_cpuid228/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid228 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid228/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid228])
        end // if (done[228])

        if (done[229]) begin
            timeout[long_cpuid229] = 0;
            //check_bad_trap(spc229_phy_pc_w, 229, long_cpuid229);
            if(active_thread[long_cpuid229])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc229_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid229/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 229 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid229]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc229_phy_pc_w))
                begin
                    if(good[long_cpuid229/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid229 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid229/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid229])
        end // if (done[229])

        if (done[230]) begin
            timeout[long_cpuid230] = 0;
            //check_bad_trap(spc230_phy_pc_w, 230, long_cpuid230);
            if(active_thread[long_cpuid230])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc230_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid230/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 230 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid230]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc230_phy_pc_w))
                begin
                    if(good[long_cpuid230/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid230 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid230/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid230])
        end // if (done[230])

        if (done[231]) begin
            timeout[long_cpuid231] = 0;
            //check_bad_trap(spc231_phy_pc_w, 231, long_cpuid231);
            if(active_thread[long_cpuid231])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc231_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid231/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 231 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid231]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc231_phy_pc_w))
                begin
                    if(good[long_cpuid231/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid231 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid231/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid231])
        end // if (done[231])

        if (done[232]) begin
            timeout[long_cpuid232] = 0;
            //check_bad_trap(spc232_phy_pc_w, 232, long_cpuid232);
            if(active_thread[long_cpuid232])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc232_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid232/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 232 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid232]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc232_phy_pc_w))
                begin
                    if(good[long_cpuid232/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid232 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid232/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid232])
        end // if (done[232])

        if (done[233]) begin
            timeout[long_cpuid233] = 0;
            //check_bad_trap(spc233_phy_pc_w, 233, long_cpuid233);
            if(active_thread[long_cpuid233])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc233_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid233/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 233 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid233]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc233_phy_pc_w))
                begin
                    if(good[long_cpuid233/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid233 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid233/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid233])
        end // if (done[233])

        if (done[234]) begin
            timeout[long_cpuid234] = 0;
            //check_bad_trap(spc234_phy_pc_w, 234, long_cpuid234);
            if(active_thread[long_cpuid234])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc234_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid234/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 234 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid234]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc234_phy_pc_w))
                begin
                    if(good[long_cpuid234/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid234 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid234/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid234])
        end // if (done[234])

        if (done[235]) begin
            timeout[long_cpuid235] = 0;
            //check_bad_trap(spc235_phy_pc_w, 235, long_cpuid235);
            if(active_thread[long_cpuid235])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc235_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid235/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 235 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid235]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc235_phy_pc_w))
                begin
                    if(good[long_cpuid235/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid235 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid235/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid235])
        end // if (done[235])

        if (done[236]) begin
            timeout[long_cpuid236] = 0;
            //check_bad_trap(spc236_phy_pc_w, 236, long_cpuid236);
            if(active_thread[long_cpuid236])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc236_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid236/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 236 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid236]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc236_phy_pc_w))
                begin
                    if(good[long_cpuid236/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid236 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid236/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid236])
        end // if (done[236])

        if (done[237]) begin
            timeout[long_cpuid237] = 0;
            //check_bad_trap(spc237_phy_pc_w, 237, long_cpuid237);
            if(active_thread[long_cpuid237])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc237_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid237/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 237 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid237]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc237_phy_pc_w))
                begin
                    if(good[long_cpuid237/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid237 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid237/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid237])
        end // if (done[237])

        if (done[238]) begin
            timeout[long_cpuid238] = 0;
            //check_bad_trap(spc238_phy_pc_w, 238, long_cpuid238);
            if(active_thread[long_cpuid238])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc238_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid238/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 238 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid238]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc238_phy_pc_w))
                begin
                    if(good[long_cpuid238/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid238 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid238/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid238])
        end // if (done[238])

        if (done[239]) begin
            timeout[long_cpuid239] = 0;
            //check_bad_trap(spc239_phy_pc_w, 239, long_cpuid239);
            if(active_thread[long_cpuid239])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc239_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid239/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 239 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid239]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc239_phy_pc_w))
                begin
                    if(good[long_cpuid239/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid239 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid239/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid239])
        end // if (done[239])

        if (done[240]) begin
            timeout[long_cpuid240] = 0;
            //check_bad_trap(spc240_phy_pc_w, 240, long_cpuid240);
            if(active_thread[long_cpuid240])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc240_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid240/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 240 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid240]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc240_phy_pc_w))
                begin
                    if(good[long_cpuid240/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid240 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid240/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid240])
        end // if (done[240])

        if (done[241]) begin
            timeout[long_cpuid241] = 0;
            //check_bad_trap(spc241_phy_pc_w, 241, long_cpuid241);
            if(active_thread[long_cpuid241])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc241_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid241/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 241 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid241]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc241_phy_pc_w))
                begin
                    if(good[long_cpuid241/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid241 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid241/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid241])
        end // if (done[241])

        if (done[242]) begin
            timeout[long_cpuid242] = 0;
            //check_bad_trap(spc242_phy_pc_w, 242, long_cpuid242);
            if(active_thread[long_cpuid242])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc242_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid242/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 242 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid242]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc242_phy_pc_w))
                begin
                    if(good[long_cpuid242/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid242 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid242/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid242])
        end // if (done[242])

        if (done[243]) begin
            timeout[long_cpuid243] = 0;
            //check_bad_trap(spc243_phy_pc_w, 243, long_cpuid243);
            if(active_thread[long_cpuid243])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc243_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid243/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 243 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid243]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc243_phy_pc_w))
                begin
                    if(good[long_cpuid243/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid243 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid243/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid243])
        end // if (done[243])

        if (done[244]) begin
            timeout[long_cpuid244] = 0;
            //check_bad_trap(spc244_phy_pc_w, 244, long_cpuid244);
            if(active_thread[long_cpuid244])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc244_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid244/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 244 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid244]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc244_phy_pc_w))
                begin
                    if(good[long_cpuid244/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid244 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid244/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid244])
        end // if (done[244])

        if (done[245]) begin
            timeout[long_cpuid245] = 0;
            //check_bad_trap(spc245_phy_pc_w, 245, long_cpuid245);
            if(active_thread[long_cpuid245])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc245_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid245/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 245 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid245]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc245_phy_pc_w))
                begin
                    if(good[long_cpuid245/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid245 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid245/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid245])
        end // if (done[245])

        if (done[246]) begin
            timeout[long_cpuid246] = 0;
            //check_bad_trap(spc246_phy_pc_w, 246, long_cpuid246);
            if(active_thread[long_cpuid246])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc246_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid246/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 246 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid246]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc246_phy_pc_w))
                begin
                    if(good[long_cpuid246/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid246 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid246/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid246])
        end // if (done[246])

        if (done[247]) begin
            timeout[long_cpuid247] = 0;
            //check_bad_trap(spc247_phy_pc_w, 247, long_cpuid247);
            if(active_thread[long_cpuid247])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc247_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid247/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 247 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid247]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc247_phy_pc_w))
                begin
                    if(good[long_cpuid247/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid247 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid247/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid247])
        end // if (done[247])

        if (done[248]) begin
            timeout[long_cpuid248] = 0;
            //check_bad_trap(spc248_phy_pc_w, 248, long_cpuid248);
            if(active_thread[long_cpuid248])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc248_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid248/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 248 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid248]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc248_phy_pc_w))
                begin
                    if(good[long_cpuid248/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid248 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid248/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid248])
        end // if (done[248])

        if (done[249]) begin
            timeout[long_cpuid249] = 0;
            //check_bad_trap(spc249_phy_pc_w, 249, long_cpuid249);
            if(active_thread[long_cpuid249])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc249_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid249/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 249 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid249]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc249_phy_pc_w))
                begin
                    if(good[long_cpuid249/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid249 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid249/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid249])
        end // if (done[249])

        if (done[250]) begin
            timeout[long_cpuid250] = 0;
            //check_bad_trap(spc250_phy_pc_w, 250, long_cpuid250);
            if(active_thread[long_cpuid250])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc250_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid250/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 250 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid250]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc250_phy_pc_w))
                begin
                    if(good[long_cpuid250/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid250 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid250/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid250])
        end // if (done[250])

        if (done[251]) begin
            timeout[long_cpuid251] = 0;
            //check_bad_trap(spc251_phy_pc_w, 251, long_cpuid251);
            if(active_thread[long_cpuid251])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc251_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid251/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 251 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid251]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc251_phy_pc_w))
                begin
                    if(good[long_cpuid251/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid251 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid251/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid251])
        end // if (done[251])

        if (done[252]) begin
            timeout[long_cpuid252] = 0;
            //check_bad_trap(spc252_phy_pc_w, 252, long_cpuid252);
            if(active_thread[long_cpuid252])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc252_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid252/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 252 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid252]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc252_phy_pc_w))
                begin
                    if(good[long_cpuid252/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid252 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid252/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid252])
        end // if (done[252])

        if (done[253]) begin
            timeout[long_cpuid253] = 0;
            //check_bad_trap(spc253_phy_pc_w, 253, long_cpuid253);
            if(active_thread[long_cpuid253])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc253_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid253/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 253 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid253]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc253_phy_pc_w))
                begin
                    if(good[long_cpuid253/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid253 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid253/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid253])
        end // if (done[253])

        if (done[254]) begin
            timeout[long_cpuid254] = 0;
            //check_bad_trap(spc254_phy_pc_w, 254, long_cpuid254);
            if(active_thread[long_cpuid254])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc254_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid254/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 254 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid254]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc254_phy_pc_w))
                begin
                    if(good[long_cpuid254/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid254 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid254/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid254])
        end // if (done[254])

        if (done[255]) begin
            timeout[long_cpuid255] = 0;
            //check_bad_trap(spc255_phy_pc_w, 255, long_cpuid255);
            if(active_thread[long_cpuid255])begin

                if(bad_trap_exists[0] & (bad_trap[0] == spc255_phy_pc_w))begin
                    hit_bad     <= 1'b1;
                    good[long_cpuid255/4]   <= 1;
                    local_diag_done = 1;
                    $display("%016t hart %4d: @@@ Hit Bad trap", $time, 255 / 4);
                    `MONITOR_PATH.fail("HIT BAD TRAP");
                end

            end
        if (active_thread[long_cpuid255]) begin
    
if(good_trap_exists[0] & (good_trap[0] == spc255_phy_pc_w))
                begin
                    if(good[long_cpuid255/4] == 0) begin
                        $display("%016t hart %4d: @@@ Hit Good trap %4d/%0d", $time, long_cpuid255 / 4, $countones(good), $bits(good));
                    end
                    good[long_cpuid255/4] <= 1'b1;
                end

            end // if (active_thread[long_cpuid255])
        end // if (done[255])

        
        end
`ifdef INCLUDE_SAS_TASKS
        get_thread_status;
`endif
        set_diag_done(local_diag_done);
    end // if (rst_l)
end // always @ (posedge clk)

always @(posedge clk) begin
  if (!rst_l) begin
    good <= '0;
    hit_bad <= 1'b0;
  end else begin
    if (&good) begin
      $display("All threads hit good tap - PASS");
      $finish;
    end
    if (hit_bad) begin
      $display("A thread hit bad trap - FAIL");
      $error;
      $finish;
    end
  end
end

endmodule


